magic
tech sky130A
magscale 1 2
timestamp 1727401017
<< nwell >>
rect -256 -819 256 819
<< pmos >>
rect -60 -600 60 600
<< pdiff >>
rect -118 588 -60 600
rect -118 -588 -106 588
rect -72 -588 -60 588
rect -118 -600 -60 -588
rect 60 588 118 600
rect 60 -588 72 588
rect 106 -588 118 588
rect 60 -600 118 -588
<< pdiffc >>
rect -106 -588 -72 588
rect 72 -588 106 588
<< nsubdiff >>
rect -220 749 -124 783
rect 124 749 220 783
rect -220 687 -186 749
rect 186 687 220 749
rect -220 -749 -186 -687
rect 186 -749 220 -687
rect -220 -783 -124 -749
rect 124 -783 220 -749
<< nsubdiffcont >>
rect -124 749 124 783
rect -220 -687 -186 687
rect 186 -687 220 687
rect -124 -783 124 -749
<< poly >>
rect -60 681 60 697
rect -60 647 -44 681
rect 44 647 60 681
rect -60 600 60 647
rect -60 -647 60 -600
rect -60 -681 -44 -647
rect 44 -681 60 -647
rect -60 -697 60 -681
<< polycont >>
rect -44 647 44 681
rect -44 -681 44 -647
<< locali >>
rect -220 749 -124 783
rect 124 749 220 783
rect -220 687 -186 749
rect 186 687 220 749
rect -60 647 -44 681
rect 44 647 60 681
rect -106 588 -72 604
rect -106 -604 -72 -588
rect 72 588 106 604
rect 72 -604 106 -588
rect -60 -681 -44 -647
rect 44 -681 60 -647
rect -220 -749 -186 -687
rect 186 -749 220 -687
rect -220 -783 -124 -749
rect 124 -783 220 -749
<< viali >>
rect -44 647 44 681
rect -106 -588 -72 588
rect 72 -588 106 588
rect -44 -681 44 -647
<< metal1 >>
rect -56 681 56 687
rect -56 647 -44 681
rect 44 647 56 681
rect -56 641 56 647
rect -112 588 -66 600
rect -112 -588 -106 588
rect -72 -588 -66 588
rect -112 -600 -66 -588
rect 66 588 112 600
rect 66 -588 72 588
rect 106 -588 112 588
rect 66 -600 112 -588
rect -56 -647 56 -641
rect -56 -681 -44 -647
rect 44 -681 56 -647
rect -56 -687 56 -681
<< properties >>
string FIXED_BBOX -203 -766 203 766
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6.0 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
