magic
tech sky130A
magscale 1 2
timestamp 1730228180
<< metal1 >>
rect 19396 31190 19596 31196
rect 19596 30990 26172 31190
rect 19396 30984 19596 30990
rect 16998 30590 17004 30790
rect 17204 30590 25772 30790
rect 14612 30190 14618 30390
rect 14818 30190 25372 30390
rect 12226 29990 12426 29996
rect 12426 29790 24976 29990
rect 12226 29784 12426 29790
rect 24776 7318 24976 29790
rect 18496 7142 24976 7318
rect 18496 7120 24776 7142
rect 18496 7118 24772 7120
rect 18496 6318 18696 7118
rect 25172 6918 25372 30190
rect 20990 6718 25372 6918
rect 20990 6318 21190 6718
rect 25572 6518 25772 30590
rect 23482 6318 25772 6518
rect 25972 6318 26172 30990
rect 17388 5913 17560 5914
rect 17388 5866 18537 5913
rect 17389 5791 18537 5866
rect 17389 2128 17575 5791
rect 30362 2800 30542 2806
rect 29848 2620 30362 2800
rect 30362 2614 30542 2620
rect 17288 2122 17676 2128
rect 17288 1728 17676 1734
rect 17276 1400 17676 1406
rect 17676 1082 18102 1318
rect 17276 994 17676 1000
rect 17882 1074 18102 1082
rect 17882 865 18553 1074
rect 17882 864 18102 865
<< via1 >>
rect 19396 30990 19596 31190
rect 17004 30590 17204 30790
rect 14618 30190 14818 30390
rect 12226 29790 12426 29990
rect 30362 2620 30542 2800
rect 17288 1734 17676 2122
rect 17276 1000 17676 1400
<< metal2 >>
rect 21862 42708 21922 42717
rect 21862 42639 21922 42648
rect 19461 42416 19470 42476
rect 19530 42416 19539 42476
rect 17078 42250 17138 42259
rect 17078 42181 17138 42190
rect 14686 42032 14746 42041
rect 14686 41963 14746 41972
rect 12294 41828 12354 41837
rect 12294 41759 12354 41768
rect 12296 41546 12352 41759
rect 14688 41584 14744 41963
rect 17080 41554 17136 42181
rect 19472 41556 19528 42416
rect 21864 41546 21920 42639
rect 12226 29990 12426 32008
rect 14618 30390 14818 32010
rect 17004 30790 17204 31992
rect 19396 31190 19596 32014
rect 21828 31642 21956 31936
rect 21828 31505 21956 31514
rect 19390 30990 19396 31190
rect 19596 30990 19602 31190
rect 17004 30584 17204 30590
rect 14618 30184 14818 30190
rect 12220 29790 12226 29990
rect 12426 29790 12432 29990
rect 30356 2620 30362 2800
rect 30542 2620 30548 2800
rect 30362 2241 30542 2620
rect 16201 2122 16579 2126
rect 16196 2117 17288 2122
rect 16196 1739 16201 2117
rect 16579 1739 17288 2117
rect 16196 1734 17288 1739
rect 17676 1734 17682 2122
rect 30358 2071 30367 2241
rect 30537 2071 30546 2241
rect 30362 2066 30542 2071
rect 16201 1730 16579 1734
rect 16181 1400 16571 1404
rect 16176 1395 17276 1400
rect 16176 1005 16181 1395
rect 16571 1005 17276 1395
rect 16176 1000 17276 1005
rect 17676 1000 17682 1400
rect 16181 996 16571 1000
<< via2 >>
rect 21862 42648 21922 42708
rect 19470 42416 19530 42476
rect 17078 42190 17138 42250
rect 14686 41972 14746 42032
rect 12294 41768 12354 41828
rect 21828 31514 21956 31642
rect 16201 1739 16579 2117
rect 30367 2071 30537 2241
rect 16181 1005 16571 1395
<< metal3 >>
rect 10320 43639 10720 43640
rect 10315 43241 10321 43639
rect 10719 43241 10725 43639
rect 27590 43628 27596 43756
rect 27724 43628 27730 43756
rect 201 42818 599 42823
rect 200 42817 1406 42818
rect 200 42419 201 42817
rect 599 42419 1406 42817
rect 200 42418 1406 42419
rect 1806 42418 1812 42818
rect 201 42413 599 42418
rect 10320 42184 10720 43241
rect 16608 42646 16614 42710
rect 16678 42708 16684 42710
rect 21857 42708 21927 42713
rect 16678 42648 21862 42708
rect 21922 42648 21927 42708
rect 16678 42646 16684 42648
rect 21857 42643 21927 42648
rect 17170 42478 17234 42484
rect 19465 42476 19535 42481
rect 17234 42416 19470 42476
rect 19530 42416 19535 42476
rect 17170 42408 17234 42414
rect 19465 42411 19535 42416
rect 17073 42250 17143 42255
rect 17718 42250 17724 42252
rect 17073 42190 17078 42250
rect 17138 42190 17724 42250
rect 17073 42185 17143 42190
rect 17718 42188 17724 42190
rect 17788 42188 17794 42252
rect 14681 42032 14751 42037
rect 18278 42034 18342 42040
rect 14681 41972 14686 42032
rect 14746 41972 18278 42032
rect 14681 41967 14751 41972
rect 18278 41964 18342 41970
rect 10320 41778 10720 41784
rect 12289 41828 12359 41833
rect 18820 41828 18826 41830
rect 12289 41768 12294 41828
rect 12354 41768 18826 41828
rect 12289 41763 12359 41768
rect 18820 41766 18826 41768
rect 18890 41766 18896 41830
rect 23054 38998 23254 39118
rect 23374 38998 23380 39118
rect 23046 34102 23294 34222
rect 23414 34102 23420 34222
rect 21823 31642 21961 31647
rect 27596 31642 27724 43628
rect 21823 31514 21828 31642
rect 21956 31514 27724 31642
rect 21823 31509 21961 31514
rect 30362 2241 30542 2246
rect 201 2128 599 2133
rect 200 2127 1392 2128
rect 200 1729 201 2127
rect 599 1729 1392 2127
rect 200 1728 1392 1729
rect 1792 1728 1798 2128
rect 14917 2127 15303 2133
rect 14916 1734 14917 2122
rect 15303 2117 16584 2122
rect 15303 1739 16201 2117
rect 16579 1739 16584 2117
rect 15303 1734 16584 1739
rect 30362 2071 30367 2241
rect 30537 2071 30542 2241
rect 201 1723 599 1728
rect 14917 1723 15303 1729
rect 14907 1400 15305 1405
rect 14906 1399 16576 1400
rect 14906 1001 14907 1399
rect 15305 1395 16576 1399
rect 15305 1005 16181 1395
rect 16571 1005 16576 1395
rect 15305 1001 16576 1005
rect 14906 1000 16576 1001
rect 14907 995 15305 1000
rect 30362 571 30542 2071
rect 30357 393 30363 571
rect 30541 393 30547 571
rect 30362 392 30542 393
<< via3 >>
rect 10321 43241 10719 43639
rect 27596 43628 27724 43756
rect 201 42419 599 42817
rect 1406 42418 1806 42818
rect 16614 42646 16678 42710
rect 17170 42414 17234 42478
rect 17724 42188 17788 42252
rect 10320 41784 10720 42184
rect 18278 41970 18342 42034
rect 18826 41766 18890 41830
rect 23254 38998 23374 39118
rect 23294 34102 23414 34222
rect 201 1729 599 2127
rect 1392 1728 1792 2128
rect 14917 1729 15303 2127
rect 14907 1001 15305 1399
rect 30363 393 30541 571
<< metal4 >>
rect 6134 44152 6194 45152
rect 6686 44152 6746 45152
rect 7238 44152 7298 45152
rect 7790 44152 7850 45152
rect 8342 44152 8402 45152
rect 8894 44152 8954 45152
rect 9446 44152 9506 45152
rect 9998 44152 10058 45152
rect 10550 44152 10610 45152
rect 11102 44152 11162 45152
rect 11654 44152 11714 45152
rect 12206 44152 12266 45152
rect 12758 44152 12818 45152
rect 13310 44152 13370 45152
rect 13862 44152 13922 45152
rect 14414 44152 14474 45152
rect 14966 44152 15026 45152
rect 15518 44152 15578 45152
rect 16070 44152 16130 45152
rect 16622 44296 16682 45152
rect 17174 44316 17234 45152
rect 16616 44170 16682 44296
rect 17172 44170 17234 44316
rect 200 42817 600 44152
rect 200 42419 201 42817
rect 599 42419 600 42817
rect 200 2127 600 42419
rect 200 1729 201 2127
rect 599 1729 600 2127
rect 200 1000 600 1729
rect 800 43752 16204 44152
rect 800 1400 1200 43752
rect 10320 43639 10720 43752
rect 10320 43241 10321 43639
rect 10719 43241 10720 43639
rect 10320 43240 10720 43241
rect 1405 42818 1807 42819
rect 1405 42418 1406 42818
rect 1806 42418 11418 42818
rect 16616 42711 16676 44170
rect 16613 42710 16679 42711
rect 16613 42646 16614 42710
rect 16678 42646 16679 42710
rect 16613 42645 16679 42646
rect 17172 42479 17232 44170
rect 1405 42417 1807 42418
rect 10319 42184 10721 42185
rect 10319 41784 10320 42184
rect 10720 41784 10721 42184
rect 10319 41783 10721 41784
rect 10320 31596 10720 41783
rect 11018 41458 11418 42418
rect 17169 42478 17235 42479
rect 17169 42414 17170 42478
rect 17234 42414 17235 42478
rect 17169 42413 17235 42414
rect 17726 42253 17786 45152
rect 18278 45000 18338 45152
rect 18272 44952 18338 45000
rect 18830 45068 18890 45152
rect 18272 44290 18332 44952
rect 18830 44796 18894 45068
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 45074 27722 45152
rect 18272 44050 18340 44290
rect 18834 44212 18894 44796
rect 17723 42252 17789 42253
rect 17723 42188 17724 42252
rect 17788 42188 17789 42252
rect 17723 42187 17789 42188
rect 18280 42035 18340 44050
rect 18828 44050 18894 44212
rect 18277 42034 18343 42035
rect 18277 41970 18278 42034
rect 18342 41970 18343 42034
rect 18277 41969 18343 41970
rect 18828 41831 18888 44050
rect 27596 43757 27724 45074
rect 28214 45050 28274 45152
rect 28766 45056 28826 45152
rect 27595 43756 27725 43757
rect 27595 43628 27596 43756
rect 27724 43628 27725 43756
rect 27595 43627 27725 43628
rect 18825 41830 18891 41831
rect 18825 41766 18826 41830
rect 18890 41766 18891 41830
rect 18825 41765 18891 41766
rect 11018 41058 21386 41458
rect 12923 39428 13243 41058
rect 15637 38340 15957 41058
rect 18351 38790 18671 41058
rect 21065 38338 21385 41058
rect 23253 39118 23375 39119
rect 28180 39118 28300 45050
rect 23253 38998 23254 39118
rect 23374 38998 28300 39118
rect 23253 38997 23375 38998
rect 23293 34222 23415 34223
rect 28760 34222 28880 45056
rect 29318 44952 29378 45152
rect 23293 34102 23294 34222
rect 23414 34102 28880 34222
rect 23293 34101 23415 34102
rect 14280 31596 14600 32588
rect 16994 31596 17314 32564
rect 19708 31596 20028 32592
rect 22422 31596 22742 32542
rect 10320 31272 22742 31596
rect 10320 31196 22740 31272
rect 1391 2128 1793 2129
rect 1391 1728 1392 2128
rect 1792 2127 15316 2128
rect 1792 1729 14917 2127
rect 15303 1729 15316 2127
rect 1792 1728 15316 1729
rect 1391 1727 1793 1728
rect 800 1399 15306 1400
rect 800 1001 14907 1399
rect 15305 1001 15306 1399
rect 800 1000 15306 1001
rect 30362 571 30542 572
rect 30362 393 30363 571
rect 30541 393 30542 571
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 393
use adc_digital_control  adc_digital_control_1
timestamp 1730221101
transform 1 0 11174 0 1 31646
box 514 0 12000 10000
use opamp_ladder  opamp_ladder_0
timestamp 1728848001
transform -1 0 28500 0 1 268
box -1708 600 10004 6050
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
