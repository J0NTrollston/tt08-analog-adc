magic
tech sky130A
magscale 1 2
timestamp 1727842972
<< metal1 >>
rect 4808 30522 4814 30722
rect 5014 30522 5828 30722
rect 18343 25802 19392 25816
rect 18343 25780 19716 25802
rect 20908 25780 20964 25786
rect 18343 25724 20908 25780
rect 18343 25703 19716 25724
rect 20908 25718 20964 25724
rect 18343 25689 19392 25703
rect 18444 19066 19214 19080
rect 18444 19040 19634 19066
rect 18444 18984 20640 19040
rect 20696 18984 20702 19040
rect 18444 18958 19634 18984
rect 18444 18944 19214 18958
rect 3478 16562 5680 16762
rect 3478 10892 3678 16562
rect 18411 12233 19184 12250
rect 18411 12206 19471 12233
rect 20392 12206 20448 12212
rect 18411 12150 20392 12206
rect 18411 12123 19471 12150
rect 20392 12144 20448 12150
rect 18411 12107 19184 12123
rect 3478 10686 3678 10692
rect 18448 5494 18914 5514
rect 18448 5472 19090 5494
rect 19472 5472 19528 5478
rect 18448 5416 19472 5472
rect 18448 5395 19090 5416
rect 19472 5410 19528 5416
rect 18448 5374 18914 5395
rect 4954 4542 4960 4742
rect 5160 4542 5724 4742
<< via1 >>
rect 4814 30522 5014 30722
rect 20908 25724 20964 25780
rect 20640 18984 20696 19040
rect 20392 12150 20448 12206
rect 3478 10692 3678 10892
rect 19472 5416 19528 5472
rect 4960 4542 5160 4742
<< metal2 >>
rect 18274 43818 18334 43827
rect 18334 43760 19924 43816
rect 18274 43749 18334 43758
rect 18832 42500 18892 42509
rect 18832 42431 18892 42440
rect 18834 41734 18890 42431
rect 19868 42178 19924 43760
rect 19868 42122 21810 42178
rect 18834 41678 19326 41734
rect 19270 39338 19326 41678
rect 21754 39416 21810 42122
rect 18718 36488 19478 36544
rect 19914 36488 20448 36544
rect 19422 36344 19478 36488
rect 19422 36288 20154 36344
rect 4814 30722 5014 30728
rect 4103 30522 4112 30722
rect 4312 30522 4814 30722
rect 4814 30516 5014 30522
rect 3472 10692 3478 10892
rect 3678 10692 3684 10892
rect 3478 2332 3678 10692
rect 20098 5472 20154 36288
rect 20392 12206 20448 36488
rect 20640 36488 21166 36544
rect 21598 36488 22362 36544
rect 20640 19040 20696 36488
rect 21598 36350 21654 36488
rect 20908 36294 21654 36350
rect 20908 25780 20964 36294
rect 20902 25724 20908 25780
rect 20964 25724 20970 25780
rect 20640 18978 20696 18984
rect 20386 12150 20392 12206
rect 20448 12150 20454 12206
rect 19466 5416 19472 5472
rect 19528 5416 20154 5472
rect 4960 4742 5160 4748
rect 4311 4542 4320 4742
rect 4520 4542 4960 4742
rect 4960 4536 5160 4542
rect 30358 2332 30558 2341
rect 3478 2132 30358 2332
rect 30358 2123 30558 2132
<< via2 >>
rect 18274 43758 18334 43818
rect 18832 42440 18892 42500
rect 4112 30522 4312 30722
rect 4320 4542 4520 4742
rect 30358 2132 30558 2332
<< metal3 >>
rect 18272 44320 18336 44326
rect 18272 44250 18336 44256
rect 18274 43823 18334 44250
rect 18269 43818 18339 43823
rect 18269 43758 18274 43818
rect 18334 43758 18339 43818
rect 18269 43753 18339 43758
rect 18830 43224 18894 43230
rect 18830 43154 18894 43160
rect 18832 42505 18892 43154
rect 18827 42500 18897 42505
rect 18827 42440 18832 42500
rect 18892 42440 18897 42500
rect 18827 42435 18897 42440
rect 19860 39253 20261 39259
rect 200 39251 18896 39252
rect 195 38853 201 39251
rect 599 38853 18896 39251
rect 200 38852 18896 38853
rect 19296 38852 19860 39252
rect 20820 39252 21220 39258
rect 20261 38852 20820 39252
rect 21220 38852 21794 39252
rect 22194 38852 22628 39252
rect 19860 38846 20261 38852
rect 20820 38846 21220 38852
rect 4107 30722 4317 30727
rect 302 30522 308 30722
rect 508 30522 4112 30722
rect 4312 30522 4317 30722
rect 4107 30517 4317 30522
rect 4315 4742 4525 4747
rect 3556 4542 3562 4742
rect 3762 4542 4320 4742
rect 4520 4542 4525 4742
rect 4315 4537 4525 4542
rect 30353 2332 30563 2337
rect 30353 2132 30358 2332
rect 30558 2132 30563 2332
rect 30353 2127 30563 2132
rect 30358 1632 30558 2127
rect 30358 1426 30558 1432
<< via3 >>
rect 18272 44256 18336 44320
rect 18830 43160 18894 43224
rect 201 38853 599 39251
rect 18896 38852 19296 39252
rect 19860 38852 20261 39253
rect 20820 38852 21220 39252
rect 21794 38852 22194 39252
rect 308 30522 508 30722
rect 3562 4542 3762 4742
rect 30358 1432 30558 1632
<< metal4 >>
rect 200 39251 600 44152
rect 200 38853 201 39251
rect 599 38853 600 39251
rect 200 30722 600 38853
rect 200 30522 308 30722
rect 508 30522 600 30722
rect 200 1000 600 30522
rect 800 43815 1200 44152
rect 6134 43815 6194 45152
rect 6686 43815 6746 45152
rect 7238 43815 7298 45152
rect 7790 43815 7850 45152
rect 8342 43815 8402 45152
rect 8894 43815 8954 45152
rect 9446 43815 9506 45152
rect 9998 43815 10058 45152
rect 10550 43815 10610 45152
rect 11102 43815 11162 45152
rect 11654 43815 11714 45152
rect 12206 43815 12266 45152
rect 12758 43815 12818 45152
rect 13310 43815 13370 45152
rect 13862 43815 13922 45152
rect 14414 43815 14474 45152
rect 14966 43815 15026 45152
rect 15518 43815 15578 45152
rect 16070 43815 16130 45152
rect 16622 43815 16682 45152
rect 17174 43815 17234 45152
rect 17726 43815 17786 45152
rect 18278 45018 18338 45152
rect 18274 44952 18338 45018
rect 18830 45032 18890 45152
rect 18830 44952 18892 45032
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 18274 44321 18334 44952
rect 18271 44320 18337 44321
rect 18271 44256 18272 44320
rect 18336 44256 18337 44320
rect 18271 44255 18337 44256
rect 800 43634 17832 43815
rect 800 39986 1200 43634
rect 18832 43225 18892 44952
rect 18829 43224 18895 43225
rect 18829 43160 18830 43224
rect 18894 43160 18895 43224
rect 18829 43159 18895 43160
rect 800 39949 22618 39986
rect 800 39586 22619 39949
rect 800 4742 1200 39586
rect 18895 39252 19297 39253
rect 18895 38852 18896 39252
rect 19296 38852 19297 39252
rect 18895 38851 19297 38852
rect 18896 38472 19296 38851
rect 19414 38392 19734 39586
rect 19859 39253 20262 39254
rect 19859 38852 19860 39253
rect 20261 38852 20262 39253
rect 19859 38851 20262 38852
rect 19897 38381 20223 38851
rect 20380 38348 20700 39586
rect 20819 39252 21221 39253
rect 20819 38852 20820 39252
rect 21220 38852 21221 39252
rect 20819 38851 21221 38852
rect 20858 38558 21182 38851
rect 21346 38392 21666 39586
rect 21793 39252 22195 39253
rect 21793 38852 21794 39252
rect 22194 38852 22195 39252
rect 21793 38851 22195 38852
rect 21832 38526 22157 38851
rect 22293 38567 22619 39586
rect 3561 4742 3763 4743
rect 800 4542 3562 4742
rect 3762 4542 3763 4742
rect 800 1000 1200 4542
rect 3561 4541 3763 4542
rect 30357 1632 30559 1633
rect 30357 1432 30358 1632
rect 30558 1432 30559 1632
rect 30357 1431 30559 1432
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30358 114 30558 1431
rect 30362 0 30542 114
use adc_digital_control  adc_digital_control_0
timestamp 1727826562
transform 1 0 18056 0 1 36488
box 514 0 4576 3000
use opamp_ladder  opamp_ladder_0
timestamp 1727841813
transform 1 0 1732 0 1 19328
box 3748 -14788 16764 11394
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
