magic
tech sky130A
magscale 1 2
timestamp 1728771870
<< error_s >>
rect 388 2115 423 2149
rect 389 2096 423 2115
rect 408 583 423 2096
rect 442 2062 477 2096
rect 847 2062 882 2079
rect 442 583 476 2062
rect 848 2061 882 2062
rect 848 2025 918 2061
rect 865 1991 936 2025
rect 1306 1991 1341 2025
rect 3770 2017 3805 2051
rect 3771 1998 3805 2017
rect 442 549 457 583
rect 865 530 935 1991
rect 1307 1972 1341 1991
rect 1783 1972 1836 1973
rect 865 494 918 530
rect 1326 477 1341 1972
rect 1360 1938 1395 1972
rect 1765 1938 1836 1972
rect 1360 477 1394 1938
rect 1766 1937 1836 1938
rect 1783 1903 1854 1937
rect 1360 443 1375 477
rect 1783 424 1853 1903
rect 2225 1284 2259 1338
rect 1783 388 1836 424
rect 2244 371 2259 1284
rect 2278 1250 2313 1284
rect 2278 371 2312 1250
rect 2424 1182 2482 1188
rect 2424 1148 2436 1182
rect 2424 1142 2482 1148
rect 2424 454 2482 460
rect 2424 420 2436 454
rect 2424 414 2482 420
rect 2278 337 2293 371
rect 2613 318 2628 1284
rect 2647 318 2681 1338
rect 3053 896 3087 914
rect 3053 860 3123 896
rect 3070 826 3141 860
rect 2647 284 2662 318
rect 3070 265 3140 826
rect 3252 758 3310 764
rect 3252 724 3264 758
rect 3252 718 3310 724
rect 3252 348 3310 354
rect 3252 314 3264 348
rect 3252 308 3310 314
rect 3070 229 3123 265
rect 3441 212 3456 860
rect 3475 212 3509 914
rect 3475 178 3490 212
rect 3790 159 3805 1998
rect 3824 1964 3859 1998
rect 4119 1964 4154 1998
rect 3824 159 3858 1964
rect 4120 1945 4154 1964
rect 3824 125 3839 159
rect 4139 106 4154 1945
rect 4173 1911 4208 1945
rect 4468 1911 4503 1945
rect 4173 106 4207 1911
rect 4469 1892 4503 1911
rect 4173 72 4188 106
rect 4488 53 4503 1892
rect 4522 1858 4557 1892
rect 4817 1858 4852 1892
rect 4522 53 4556 1858
rect 4818 1839 4852 1858
rect 4522 19 4537 53
rect 4837 0 4852 1839
rect 4871 1805 4906 1839
rect 4871 0 4905 1805
rect 4871 -34 4886 0
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use sky130_fd_pr__pfet_01v8_XPP7BA  XM1
timestamp 1728771870
transform 1 0 203 0 1 1366
box -256 -819 256 819
use sky130_fd_pr__pfet_01v8_XPP7BA  XM2
timestamp 1728771870
transform 1 0 662 0 1 1313
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_3BHWKV  XM3
timestamp 1728771870
transform 1 0 1121 0 1 1251
box -256 -810 256 810
use sky130_fd_pr__nfet_01v8_3BHWKV  XM4
timestamp 1728771870
transform 1 0 1580 0 1 1198
box -256 -810 256 810
use sky130_fd_pr__pfet_01v8_XPP7BA  XM5
timestamp 1728771870
transform 1 0 2039 0 1 1154
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_848SAM  XM6
timestamp 1728771870
transform 1 0 3281 0 1 536
box -211 -360 211 360
use sky130_fd_pr__pfet_01v8_XGSNAL  XM7
timestamp 1728771870
transform 1 0 2453 0 1 801
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XPP7BA  XM8
timestamp 1728771870
transform 1 0 2867 0 1 1048
box -256 -819 256 819
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR1
timestamp 1728771870
transform 1 0 3989 0 1 1052
box -201 -982 201 982
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR2
timestamp 1728771870
transform 1 0 4338 0 1 999
box -201 -982 201 982
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR3
timestamp 1728771870
transform 1 0 4687 0 1 946
box -201 -982 201 982
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR4
timestamp 1728771870
transform 1 0 5036 0 1 893
box -201 -982 201 982
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR
timestamp 1728771870
transform 1 0 3640 0 1 1105
box -201 -982 201 982
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 vin_n
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 vin_p
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vout
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VGND
port 4 nsew
<< end >>
