magic
tech sky130A
magscale 1 2
timestamp 1727813169
<< pwell >>
rect -258 -1101 258 1101
<< ndiff >>
rect -100 931 100 943
rect -100 897 -88 931
rect 88 897 100 931
rect -100 840 100 897
rect -100 -897 100 -840
rect -100 -931 -88 -897
rect 88 -931 100 -897
rect -100 -943 100 -931
<< ndiffc >>
rect -88 897 88 931
rect -88 -931 88 -897
<< psubdiff >>
rect -222 1031 -126 1065
rect 126 1031 222 1065
rect -222 969 -188 1031
rect 188 969 222 1031
rect -222 -1031 -188 -969
rect 188 -1031 222 -969
rect -222 -1065 -126 -1031
rect 126 -1065 222 -1031
<< psubdiffcont >>
rect -126 1031 126 1065
rect -222 -969 -188 969
rect 188 -969 222 969
rect -126 -1065 126 -1031
<< ndiffres >>
rect -100 -840 100 840
<< locali >>
rect -222 1031 -126 1065
rect 126 1031 222 1065
rect -222 969 -188 1031
rect 188 969 222 1031
rect -104 897 -88 931
rect 88 897 104 931
rect -104 -931 -88 -897
rect 88 -931 104 -897
rect -222 -1031 -188 -969
rect 188 -1031 222 -969
rect -222 -1065 -126 -1031
rect 126 -1065 222 -1031
<< viali >>
rect -88 897 88 931
rect -88 857 88 897
rect -88 -897 88 -857
rect -88 -931 88 -897
<< metal1 >>
rect -100 931 100 937
rect -100 857 -88 931
rect 88 857 100 931
rect -100 851 100 857
rect -100 -857 100 -851
rect -100 -931 -88 -857
rect 88 -931 100 -857
rect -100 -937 100 -931
<< properties >>
string FIXED_BBOX -205 -1048 205 1048
string gencell sky130_fd_pr__res_generic_nd
string library sky130
string parameters w 1.0 l 8.4 m 1 nx 1 wmin 0.42 lmin 2.10 rho 120 val 1.061k dummy 0 dw 0.05 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
