magic
tech sky130A
magscale 1 2
timestamp 1728800409
<< pwell >>
rect 8840 1146 8888 1346
rect 8910 -740 9016 -494
<< viali >>
rect 7754 3522 9004 3556
rect 6880 1238 6914 1468
rect 6968 1272 7002 1468
rect 6968 1238 7298 1272
rect 7352 1238 7682 1272
rect 6968 1132 7298 1166
rect 6968 -726 7298 -692
rect 7352 -1022 7386 -692
rect 7352 -1162 7682 -1128
rect 7754 -1162 8600 -1128
rect 8654 -1162 9004 -1128
<< metal1 >>
rect 6548 3556 9040 3722
rect 6548 3522 7754 3556
rect 9004 3522 9040 3556
rect 7718 3516 9040 3522
rect 8058 3374 8296 3516
rect 8654 3374 8768 3516
rect 8796 3414 8862 3470
rect 7718 3000 7902 3374
rect 6714 2568 7168 3000
rect 7482 2568 7902 3000
rect 7718 2208 7902 2568
rect 7718 2132 7908 2208
rect 8046 2172 8308 3374
rect 8452 2172 8544 3374
rect 8654 2772 8802 3374
rect 8850 2772 9040 3374
rect 7718 2076 8440 2132
rect 8498 2036 8544 2172
rect 8148 1978 8544 2036
rect 8666 2676 8862 2732
rect 8148 1842 8206 1978
rect 6874 1468 7026 1480
rect 6714 1036 6784 1396
rect 6874 1238 6880 1468
rect 6914 1238 6968 1468
rect 7002 1278 7026 1468
rect 7098 1368 7552 1800
rect 7002 1272 7694 1278
rect 7298 1238 7352 1272
rect 7682 1238 7694 1272
rect 6874 1166 7694 1238
rect 6874 1132 6968 1166
rect 7298 1132 7694 1166
rect 6874 1126 7694 1132
rect 6714 604 7168 1036
rect 7822 640 7902 1842
rect 8040 640 8314 1842
rect 8446 1832 8550 1842
rect 8452 640 8550 1832
rect 6802 520 6890 526
rect 6548 346 6748 402
rect 6802 346 6890 432
rect 6548 258 6890 346
rect 6548 202 6748 258
rect 7280 168 7552 600
rect 7822 300 7890 640
rect 7930 520 8018 594
rect 7930 426 8018 432
rect 8336 520 8424 594
rect 8336 426 8424 432
rect 8470 490 8550 640
rect 8666 490 8796 2676
rect 8910 1346 9040 2772
rect 8840 1146 9040 1346
rect 8470 354 8796 490
rect 7822 244 8440 300
rect 7822 212 7890 244
rect 8470 212 8550 354
rect 6548 -58 6748 2
rect 6548 -146 6800 -58
rect 6888 -146 6894 -58
rect 6548 -198 6748 -146
rect 7280 -164 7352 168
rect 7098 -596 7352 -164
rect 7346 -686 7392 -680
rect 6956 -692 7392 -686
rect 6956 -726 6968 -692
rect 7298 -726 7352 -692
rect 6956 -732 7352 -726
rect 7346 -1022 7352 -732
rect 7386 -1022 7392 -692
rect 7822 -988 7902 212
rect 8046 -988 8308 212
rect 8452 -982 8550 212
rect 8666 -600 8796 354
rect 8666 -656 8862 -600
rect 8910 -688 9040 1146
rect 8452 -988 8466 -982
rect 7346 -1034 7392 -1022
rect 7482 -1122 7552 -1002
rect 8058 -1122 8296 -988
rect 8470 -994 8550 -982
rect 8654 -988 8802 -688
rect 8856 -988 9040 -688
rect 8654 -1122 8768 -988
rect 8796 -1076 8862 -1020
rect 7340 -1128 9040 -1122
rect 6548 -1162 7352 -1128
rect 7682 -1162 7754 -1128
rect 8600 -1162 8654 -1128
rect 9004 -1162 9040 -1128
rect 6548 -1328 9040 -1162
<< via1 >>
rect 6802 432 6890 520
rect 7930 432 8018 520
rect 8336 432 8424 520
rect 6800 -146 6888 -58
<< metal2 >>
rect 8326 520 8434 530
rect 6796 432 6802 520
rect 6890 432 7930 520
rect 8018 432 8024 520
rect 8326 432 8336 520
rect 8424 432 8434 520
rect 8326 422 8434 432
rect 6805 144 6883 148
rect 6800 139 6888 144
rect 6800 61 6805 139
rect 6883 61 6888 139
rect 6800 -58 6888 61
rect 6800 -152 6888 -146
<< via2 >>
rect 8336 432 8424 520
rect 6805 61 6883 139
<< metal3 >>
rect 8331 520 8429 525
rect 8132 432 8336 520
rect 8424 432 8429 520
rect 8132 414 8220 432
rect 8331 427 8429 432
rect 8336 422 8424 427
rect 6988 326 8220 414
rect 6988 144 7076 326
rect 6800 139 7076 144
rect 6800 61 6805 139
rect 6883 61 7076 139
rect 6800 56 7076 61
use sky130_fd_pr__pfet_01v8_XPP7BA  XM1
timestamp 1728771870
transform 1 0 7974 0 1 1241
box -256 -819 256 819
use sky130_fd_pr__pfet_01v8_XPP7BA  XM2
timestamp 1728771870
transform 1 0 8380 0 1 1241
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_3BHWKV  XM3
timestamp 1728771870
transform 1 0 7974 0 1 -388
box -256 -810 256 810
use sky130_fd_pr__nfet_01v8_3BHWKV  XM4
timestamp 1728771870
transform 1 0 8380 0 1 -388
box -256 -810 256 810
use sky130_fd_pr__pfet_01v8_XPP7BA  XM5
timestamp 1728771870
transform 1 0 8380 0 1 2773
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_848SAM  XM6
timestamp 1728771870
transform 1 0 8829 0 1 -838
box -211 -360 211 360
use sky130_fd_pr__pfet_01v8_XGSNAL  XM7
timestamp 1728771870
transform 1 0 8829 0 1 3073
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XPP7BA  XM8
timestamp 1728771870
transform 1 0 7974 0 1 2773
box -256 -819 256 819
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR1
timestamp 1728771870
transform 1 0 7133 0 1 220
box -201 -982 201 982
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR2
timestamp 1728771870
transform 1 0 6749 0 1 2184
box -201 -982 201 982
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR3
timestamp 1728771870
transform 1 0 7133 0 1 2184
box -201 -982 201 982
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR4
timestamp 1728771870
transform 1 0 7517 0 1 2184
box -201 -982 201 982
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR
timestamp 1728771870
transform 1 0 7517 0 1 -216
box -201 -982 201 982
<< labels >>
flabel metal1 8840 1146 9040 1346 0 FreeSans 256 0 0 0 Vout
port 3 nsew
flabel metal1 6548 3522 6748 3722 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 6548 -1328 6748 -1128 0 FreeSans 256 0 0 0 VGND
port 4 nsew
flabel metal1 6548 202 6748 402 0 FreeSans 256 0 0 0 vin_n
port 1 nsew
flabel metal1 6548 -198 6748 2 0 FreeSans 256 0 0 0 vin_p
port 2 nsew
<< end >>
