magic
tech sky130A
magscale 1 2
timestamp 1728849390
<< metal1 >>
rect 25966 39788 25972 39988
rect 26172 39788 26178 39988
rect 25572 39588 25772 39594
rect 25172 39188 25372 39194
rect 24772 38788 24972 38794
rect 24772 7318 24972 38588
rect 18496 7118 24972 7318
rect 18496 6318 18696 7118
rect 25172 6918 25372 38988
rect 20990 6718 25372 6918
rect 20990 6318 21190 6718
rect 25572 6518 25772 39388
rect 23482 6318 25772 6518
rect 25972 6318 26172 39788
rect 17388 5913 17560 5914
rect 17388 5866 18537 5913
rect 17389 5791 18537 5866
rect 17389 2128 17575 5791
rect 30362 2800 30542 2806
rect 29848 2620 30362 2800
rect 30362 2614 30542 2620
rect 17288 2122 17676 2128
rect 17288 1728 17676 1734
rect 17276 1400 17676 1406
rect 17676 1082 18102 1318
rect 17276 994 17676 1000
rect 17882 1074 18102 1082
rect 17882 865 18553 1074
rect 17882 864 18102 865
<< via1 >>
rect 25972 39788 26172 39988
rect 25572 39388 25772 39588
rect 25172 38988 25372 39188
rect 24772 38588 24972 38788
rect 30362 2620 30542 2800
rect 17288 1734 17676 2122
rect 17276 1000 17676 1400
<< metal2 >>
rect 18834 42894 18894 42903
rect 18294 42836 18834 42892
rect 18834 42825 18894 42834
rect 19122 42894 19182 42903
rect 19182 42836 20834 42892
rect 19122 42825 19182 42834
rect 17670 38788 17870 39992
rect 18866 39188 19066 39990
rect 25972 39988 26172 39994
rect 20062 39588 20262 39988
rect 21260 39788 25972 39988
rect 25972 39782 26172 39788
rect 20062 39388 25572 39588
rect 25772 39388 25778 39588
rect 18866 38988 25172 39188
rect 25372 38988 25378 39188
rect 17670 38588 24772 38788
rect 24972 38588 24978 38788
rect 30356 2620 30362 2800
rect 30542 2620 30548 2800
rect 30362 2241 30542 2620
rect 16201 2122 16579 2126
rect 16196 2117 17288 2122
rect 16196 1739 16201 2117
rect 16579 1739 17288 2117
rect 16196 1734 17288 1739
rect 17676 1734 17682 2122
rect 30358 2071 30367 2241
rect 30537 2071 30546 2241
rect 30362 2066 30542 2071
rect 16201 1730 16579 1734
rect 16181 1400 16571 1404
rect 16176 1395 17276 1400
rect 16176 1005 16181 1395
rect 16571 1005 17276 1395
rect 16176 1000 17276 1005
rect 17676 1000 17682 1400
rect 16181 996 16571 1000
<< via2 >>
rect 18834 42834 18894 42894
rect 19122 42834 19182 42894
rect 16201 1739 16579 2117
rect 30367 2071 30537 2241
rect 16181 1005 16571 1395
<< metal3 >>
rect 18832 43780 18896 43786
rect 18832 43710 18896 43716
rect 16770 43613 17170 43614
rect 16765 43215 16771 43613
rect 17169 43215 17175 43613
rect 201 42818 599 42823
rect 200 42817 1406 42818
rect 200 42419 201 42817
rect 599 42419 1406 42817
rect 200 42418 1406 42419
rect 1806 42418 1812 42818
rect 201 42413 599 42418
rect 16770 42088 17170 43215
rect 18834 42899 18894 43710
rect 19120 43338 19184 43344
rect 19120 43268 19184 43274
rect 19122 42899 19182 43268
rect 18829 42894 18899 42899
rect 18829 42834 18834 42894
rect 18894 42834 18899 42894
rect 18829 42829 18899 42834
rect 19117 42894 19187 42899
rect 19117 42834 19122 42894
rect 19182 42834 19187 42894
rect 19117 42829 19187 42834
rect 16770 41682 17170 41688
rect 30362 2241 30542 2246
rect 201 2128 599 2133
rect 200 2127 1392 2128
rect 200 1729 201 2127
rect 599 1729 1392 2127
rect 200 1728 1392 1729
rect 1792 1728 1798 2128
rect 14917 2127 15303 2133
rect 14916 1734 14917 2122
rect 15303 2117 16584 2122
rect 15303 1739 16201 2117
rect 16579 1739 16584 2117
rect 15303 1734 16584 1739
rect 30362 2071 30367 2241
rect 30537 2071 30542 2241
rect 201 1723 599 1728
rect 14917 1723 15303 1729
rect 14907 1400 15305 1405
rect 14906 1399 16576 1400
rect 14906 1001 14907 1399
rect 15305 1395 16576 1399
rect 15305 1005 16181 1395
rect 16571 1005 16576 1395
rect 15305 1001 16576 1005
rect 14906 1000 16576 1001
rect 14907 995 15305 1000
rect 30362 571 30542 2071
rect 30357 393 30363 571
rect 30541 393 30547 571
rect 30362 392 30542 393
<< via3 >>
rect 18832 43716 18896 43780
rect 16771 43215 17169 43613
rect 201 42419 599 42817
rect 1406 42418 1806 42818
rect 19120 43274 19184 43338
rect 16770 41688 17170 42088
rect 201 1729 599 2127
rect 1392 1728 1792 2128
rect 14917 1729 15303 2127
rect 14907 1001 15305 1399
rect 30363 393 30541 571
<< metal4 >>
rect 6134 44152 6194 45152
rect 6686 44152 6746 45152
rect 7238 44152 7298 45152
rect 7790 44152 7850 45152
rect 8342 44152 8402 45152
rect 8894 44152 8954 45152
rect 9446 44152 9506 45152
rect 9998 44152 10058 45152
rect 10550 44152 10610 45152
rect 11102 44152 11162 45152
rect 11654 44152 11714 45152
rect 12206 44152 12266 45152
rect 12758 44152 12818 45152
rect 13310 44152 13370 45152
rect 13862 44152 13922 45152
rect 14414 44152 14474 45152
rect 14966 44152 15026 45152
rect 15518 44152 15578 45152
rect 16070 44152 16130 45152
rect 16622 44152 16682 45152
rect 17174 44152 17234 45152
rect 17726 44152 17786 45152
rect 18278 45000 18338 45152
rect 18272 44952 18338 45000
rect 18830 45068 18890 45152
rect 200 42817 600 44152
rect 200 42419 201 42817
rect 599 42419 600 42817
rect 200 2127 600 42419
rect 200 1729 201 2127
rect 599 1729 600 2127
rect 200 1000 600 1729
rect 800 43752 17828 44152
rect 800 1400 1200 43752
rect 16770 43613 17170 43752
rect 16770 43215 16771 43613
rect 17169 43215 17170 43613
rect 18272 43336 18332 44952
rect 18830 44796 18894 45068
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 18834 43781 18894 44796
rect 18831 43780 18897 43781
rect 18831 43716 18832 43780
rect 18896 43716 18897 43780
rect 18831 43715 18897 43716
rect 19119 43338 19185 43339
rect 19119 43336 19120 43338
rect 18272 43276 19120 43336
rect 19119 43274 19120 43276
rect 19184 43274 19185 43338
rect 19119 43273 19185 43274
rect 16770 43214 17170 43215
rect 1405 42818 1807 42819
rect 1405 42418 1406 42818
rect 1806 42418 21173 42818
rect 1405 42417 1807 42418
rect 16769 42088 17171 42089
rect 16769 41688 16770 42088
rect 17170 41688 17171 42088
rect 16769 41687 17171 41688
rect 16770 40034 17170 41687
rect 17955 41598 18275 42418
rect 18921 41564 19241 42418
rect 19887 41588 20207 42418
rect 20853 41518 21173 42418
rect 18438 40034 18758 41492
rect 19404 40034 19724 40788
rect 20370 40034 20690 40792
rect 21336 40034 21656 40788
rect 16770 39634 21656 40034
rect 1391 2128 1793 2129
rect 1391 1728 1392 2128
rect 1792 2127 15316 2128
rect 1792 1729 14917 2127
rect 15303 1729 15316 2127
rect 1792 1728 15316 1729
rect 1391 1727 1793 1728
rect 800 1399 15306 1400
rect 800 1001 14907 1399
rect 15305 1001 15306 1399
rect 800 1000 15306 1001
rect 30362 571 30542 572
rect 30362 393 30363 571
rect 30541 393 30542 571
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 393
use adc_digital_control  adc_digital_control_0
timestamp 1727826562
transform 1 0 17080 0 1 39892
box 514 0 4576 3000
use opamp_ladder  opamp_ladder_0
timestamp 1728848001
transform -1 0 28500 0 1 268
box -1708 600 10004 6050
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
