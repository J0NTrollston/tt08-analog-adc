magic
tech sky130A
magscale 1 2
timestamp 1728450646
<< nwell >>
rect 18902 42223 19223 42882
<< metal1 >>
rect 18660 33872 19220 33878
rect 17472 33796 18032 33802
rect 17472 26072 18032 33236
rect 21054 33872 21614 33878
rect 18660 26088 19220 33312
rect 19858 33796 20418 33802
rect 19858 26194 20418 33236
rect 21054 26194 21614 33312
rect 19852 25634 19858 26194
rect 20418 25634 20424 26194
rect 21048 25634 21054 26194
rect 21614 25634 21620 26194
rect 18660 25522 19220 25528
rect 17472 25506 18032 25512
rect 17466 21908 18026 21914
rect 17466 20270 18026 21348
rect 13474 20230 14034 20236
rect 17466 19704 18026 19710
rect 13474 19042 14034 19670
rect 13468 18482 13474 19042
rect 14034 18482 14040 19042
rect 18654 18986 18660 19546
rect 19220 18986 19226 19546
rect 8162 17940 8722 17946
rect 8162 16116 8722 17380
rect 15868 16688 15874 17248
rect 16434 16688 16440 17248
rect 18660 17208 19220 18986
rect 8156 15556 8162 16116
rect 8722 15556 8728 16116
rect 15874 15660 16434 16688
rect 18660 16642 19220 16648
rect 15874 15094 16434 15100
rect 3872 4036 4272 4042
rect 4272 3636 29582 3640
rect 3872 3240 29582 3636
rect 2323 3111 2725 3117
rect 2725 2709 3529 3111
rect 2323 2703 2725 2709
rect 17239 767 17521 1499
rect 17233 485 17239 767
rect 17521 485 17527 767
<< via1 >>
rect 17472 33236 18032 33796
rect 17472 25512 18032 26072
rect 18660 33312 19220 33872
rect 19858 33236 20418 33796
rect 21054 33312 21614 33872
rect 18660 25528 19220 26088
rect 19858 25634 20418 26194
rect 21054 25634 21614 26194
rect 17466 21348 18026 21908
rect 13474 19670 14034 20230
rect 17466 19710 18026 20270
rect 13474 18482 14034 19042
rect 18660 18986 19220 19546
rect 8162 17380 8722 17940
rect 15874 16688 16434 17248
rect 8162 15556 8722 16116
rect 18660 16648 19220 17208
rect 15874 15100 16434 15660
rect 3872 3636 4272 4036
rect 2323 2709 2725 3111
rect 17239 485 17521 767
<< metal2 >>
rect 19774 43666 19783 43773
rect 19890 43666 20842 43773
rect 18247 43631 18362 43640
rect 18247 43237 18362 43516
rect 20735 43243 20842 43666
rect 21326 40739 21354 40774
rect 17676 40548 17829 40704
rect 17598 39712 17907 40548
rect 18861 40543 19019 40731
rect 20058 40559 20218 40722
rect 21259 40575 21409 40739
rect 17472 33796 18032 39712
rect 18779 39704 19101 40543
rect 19973 39712 20303 40559
rect 21175 39720 21493 40575
rect 18660 33872 19220 39704
rect 17466 33236 17472 33796
rect 18032 33236 18038 33796
rect 18654 33312 18660 33872
rect 19220 33312 19226 33872
rect 19858 33796 20418 39712
rect 21054 33872 21614 39720
rect 19852 33236 19858 33796
rect 20418 33236 20424 33796
rect 21048 33312 21054 33872
rect 21614 33312 21620 33872
rect 19858 26194 20418 26200
rect 17466 25512 17472 26072
rect 18032 25512 18038 26072
rect 18654 25528 18660 26088
rect 19220 25528 19226 26088
rect 17472 24046 18032 25512
rect 17466 23678 18032 24046
rect 17466 21908 18026 23678
rect 17460 21348 17466 21908
rect 18026 21348 18032 21908
rect 13468 19670 13474 20230
rect 14034 19670 14632 20230
rect 15192 19670 15201 20230
rect 16607 19710 16616 20270
rect 17176 19710 17466 20270
rect 18026 19710 18032 20270
rect 18660 19546 19220 25528
rect 19858 19575 20418 25634
rect 21054 26194 21614 26200
rect 21054 19651 21614 25634
rect 13474 19042 14034 19048
rect 19854 19025 19863 19575
rect 20413 19025 20422 19575
rect 21050 19101 21059 19651
rect 21609 19101 21618 19651
rect 21054 19096 21614 19101
rect 19858 19020 20418 19025
rect 18660 18980 19220 18986
rect 8156 17380 8162 17940
rect 8722 17380 9618 17940
rect 10178 17380 10187 17940
rect 13474 17935 14034 18482
rect 21054 18395 21614 18400
rect 13474 17385 13479 17935
rect 14029 17385 14034 17935
rect 21050 17845 21059 18395
rect 21609 17845 21618 18395
rect 13474 17380 14034 17385
rect 19858 17775 20413 17784
rect 13479 17376 14029 17380
rect 15874 17248 16434 17254
rect 16434 17208 18392 17248
rect 16434 16688 18660 17208
rect 15874 16682 16434 16688
rect 17892 16648 18660 16688
rect 19220 16648 19226 17208
rect 6706 16116 7266 16134
rect 8162 16116 8722 16122
rect 6706 15556 8162 16116
rect 19858 16012 20413 17220
rect 6706 15021 7266 15556
rect 8162 15550 8722 15556
rect 6706 14471 6711 15021
rect 7261 14471 7266 15021
rect 13502 15155 15874 15660
rect 13502 14605 13507 15155
rect 14057 15100 15874 15155
rect 16434 15100 16440 15660
rect 21054 16092 21614 17845
rect 24839 15734 25389 15738
rect 21054 15523 21614 15532
rect 19858 15448 20413 15457
rect 22385 15174 22394 15734
rect 22954 15729 25394 15734
rect 22954 15179 24839 15729
rect 25389 15179 25394 15729
rect 22954 15174 25394 15179
rect 24839 15170 25389 15174
rect 14057 14605 14062 15100
rect 13502 14600 14062 14605
rect 13507 14596 14057 14600
rect 6706 14466 7266 14471
rect 6711 14462 7261 14466
rect 2197 4036 2587 4040
rect 2192 4031 3872 4036
rect 2192 3641 2197 4031
rect 2587 3641 3872 4031
rect 2192 3636 3872 3641
rect 4272 3636 4278 4036
rect 2197 3632 2587 3636
rect 1666 3111 2058 3115
rect 1661 3106 2323 3111
rect 1661 2714 1666 3106
rect 2058 2714 2323 3106
rect 1661 2709 2323 2714
rect 2725 2709 2731 3111
rect 1666 2705 2058 2709
rect 17239 767 17521 773
rect 18772 767 19044 771
rect 17521 762 19049 767
rect 17521 490 18772 762
rect 19044 490 19049 762
rect 17521 485 19049 490
rect 17239 479 17521 485
rect 18772 481 19044 485
<< via2 >>
rect 19783 43666 19890 43773
rect 18247 43516 18362 43631
rect 14632 19670 15192 20230
rect 16616 19710 17176 20270
rect 19863 19025 20413 19575
rect 21059 19101 21609 19651
rect 9618 17380 10178 17940
rect 13479 17385 14029 17935
rect 21059 17845 21609 18395
rect 19858 17220 20413 17775
rect 6711 14471 7261 15021
rect 13507 14605 14057 15155
rect 19858 15457 20413 16012
rect 21054 15532 21614 16092
rect 22394 15174 22954 15734
rect 24839 15179 25389 15729
rect 2197 3641 2587 4031
rect 1666 2714 2058 3106
rect 18772 490 19044 762
<< metal3 >>
rect 18241 43900 18247 44015
rect 18362 43900 18368 44015
rect 16730 43814 17131 43815
rect 16722 43415 16728 43814
rect 17133 43415 17139 43814
rect 18247 43636 18362 43900
rect 19778 43773 19895 43778
rect 18797 43666 18803 43773
rect 18910 43666 19783 43773
rect 19890 43666 19895 43773
rect 19778 43661 19895 43666
rect 18242 43631 18367 43636
rect 18242 43516 18247 43631
rect 18362 43516 18367 43631
rect 18242 43511 18367 43516
rect 1952 43090 2352 43096
rect 196 42690 202 43090
rect 602 42690 1952 43090
rect 1952 42684 2352 42690
rect 16730 40595 17131 43415
rect 16730 40188 17131 40194
rect 16611 20270 17181 20275
rect 14627 20230 15197 20235
rect 15594 20230 16616 20270
rect 14627 19670 14632 20230
rect 15192 19710 16616 20230
rect 17176 19710 17181 20270
rect 15192 19670 15738 19710
rect 16611 19705 17181 19710
rect 14627 19665 15197 19670
rect 21054 19651 21614 19656
rect 19858 19575 20418 19580
rect 19858 19025 19863 19575
rect 20413 19025 20418 19575
rect 19858 18470 20418 19025
rect 21054 19101 21059 19651
rect 21609 19101 21614 19651
rect 9613 17940 10183 17945
rect 12113 17940 12671 17945
rect 9613 17380 9618 17940
rect 10178 17380 10850 17940
rect 11410 17380 11416 17940
rect 12112 17939 14034 17940
rect 12112 17381 12113 17939
rect 12671 17935 14034 17939
rect 12671 17385 13479 17935
rect 14029 17385 14034 17935
rect 19858 17780 20413 18470
rect 21054 18395 21614 19101
rect 21054 17845 21059 18395
rect 21609 17845 21614 18395
rect 21054 17840 21614 17845
rect 12671 17381 14034 17385
rect 12112 17380 14034 17381
rect 19853 17775 20418 17780
rect 9613 17375 10183 17380
rect 12113 17375 12671 17380
rect 19853 17220 19858 17775
rect 20413 17220 20418 17775
rect 19853 17215 20418 17220
rect 19858 16017 20418 16100
rect 21054 16097 21614 16100
rect 19853 16012 20418 16017
rect 19853 15722 19858 16012
rect 19370 15654 19858 15722
rect 19064 15457 19858 15654
rect 20413 15457 20418 16012
rect 21049 16092 21619 16097
rect 21049 15532 21054 16092
rect 21614 15734 21619 16092
rect 22389 15734 22959 15739
rect 21614 15532 22394 15734
rect 21049 15527 22394 15532
rect 19064 15162 20418 15457
rect 21054 15174 22394 15527
rect 22954 15174 22959 15734
rect 24834 15729 26400 15734
rect 24834 15179 24839 15729
rect 25389 15179 26400 15729
rect 24834 15174 26400 15179
rect 22389 15169 22959 15174
rect 12246 15155 14062 15160
rect 5522 15021 7266 15026
rect 5522 14471 6711 15021
rect 7261 14471 7266 15021
rect 5522 14466 7266 14471
rect 12246 14605 13507 15155
rect 14057 14605 14062 15155
rect 12246 14600 14062 14605
rect 5522 14341 6082 14466
rect 12246 14461 12806 14600
rect 19064 14533 19624 15162
rect 25840 14539 26400 15174
rect 5522 13783 5523 14341
rect 6081 13783 6082 14341
rect 12241 13903 12247 14461
rect 12805 13903 12811 14461
rect 19059 13975 19065 14533
rect 19623 13975 19629 14533
rect 25835 13981 25841 14539
rect 26399 13981 26405 14539
rect 25840 13980 26400 13981
rect 19064 13974 19624 13975
rect 12246 13902 12806 13903
rect 5522 13782 6082 13783
rect 5523 13777 6081 13782
rect 1459 4036 1857 4041
rect 1458 4035 2592 4036
rect 1458 3637 1459 4035
rect 1857 4031 2592 4035
rect 1857 3641 2197 4031
rect 2587 3641 2592 4031
rect 1857 3637 2592 3641
rect 1458 3636 2592 3637
rect 1459 3631 1857 3636
rect 201 3110 599 3115
rect 1447 3110 2063 3111
rect 200 3109 2063 3110
rect 200 2711 201 3109
rect 599 3106 2063 3109
rect 599 2714 1666 3106
rect 2058 2714 2063 3106
rect 599 2711 2063 2714
rect 200 2710 2063 2711
rect 201 2705 599 2710
rect 1447 2709 2063 2710
rect 19542 767 19844 776
rect 18767 766 19844 767
rect 18767 762 19552 766
rect 18767 490 18772 762
rect 19044 490 19552 762
rect 18767 486 19552 490
rect 19832 486 19844 766
rect 18767 485 19844 486
rect 19542 474 19844 485
<< via3 >>
rect 18247 43900 18362 44015
rect 16728 43415 17133 43814
rect 18803 43666 18910 43773
rect 202 42690 602 43090
rect 1952 42690 2352 43090
rect 16730 40194 17131 40595
rect 10850 17380 11410 17940
rect 12113 17381 12671 17939
rect 5523 13783 6081 14341
rect 12247 13903 12805 14461
rect 19065 13975 19623 14533
rect 25841 13981 26399 14539
rect 1459 3637 1857 4035
rect 201 2711 599 3109
rect 19552 486 19832 766
<< metal4 >>
rect 200 43091 600 44152
rect 800 43815 1200 44152
rect 6134 43815 6194 45152
rect 6686 43815 6746 45152
rect 7238 43815 7298 45152
rect 7790 43815 7850 45152
rect 8342 43815 8402 45152
rect 8894 43815 8954 45152
rect 9446 43815 9506 45152
rect 9998 43815 10058 45152
rect 10550 43815 10610 45152
rect 11102 43815 11162 45152
rect 11654 43815 11714 45152
rect 12206 43815 12266 45152
rect 12758 43815 12818 45152
rect 13310 43815 13370 45152
rect 13862 43815 13922 45152
rect 14414 43815 14474 45152
rect 14966 43815 15026 45152
rect 15518 43815 15578 45152
rect 16070 43815 16130 45152
rect 16622 43815 16682 45152
rect 17174 43815 17234 45152
rect 17726 43815 17786 45152
rect 18278 45018 18338 45152
rect 18274 44952 18338 45018
rect 18830 45032 18890 45152
rect 18830 44952 18892 45032
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 18274 44841 18334 44952
rect 18832 44843 18892 44952
rect 18241 44015 18367 44841
rect 18241 43900 18247 44015
rect 18362 43900 18367 44015
rect 18241 43894 18367 43900
rect 800 43814 17834 43815
rect 800 43415 16728 43814
rect 17133 43415 17834 43814
rect 18803 43774 18910 44843
rect 18802 43773 18911 43774
rect 18802 43666 18803 43773
rect 18910 43666 18911 43773
rect 18802 43665 18911 43666
rect 800 43414 17834 43415
rect 200 43090 603 43091
rect 200 42690 202 43090
rect 602 42690 603 43090
rect 200 42689 603 42690
rect 200 3109 600 42689
rect 200 2711 201 3109
rect 599 2711 600 3109
rect 200 1000 600 2711
rect 800 4036 1200 43414
rect 1951 43090 2353 43091
rect 20835 43090 21155 43094
rect 1951 42690 1952 43090
rect 2352 42690 21155 43090
rect 1951 42689 2353 42690
rect 17937 41996 18257 42690
rect 19869 42154 20189 42690
rect 20835 42154 21155 42690
rect 16729 40595 17132 40596
rect 17454 40595 17774 41226
rect 18420 40595 18740 41322
rect 19386 40595 19706 41226
rect 20352 40595 20672 41226
rect 16729 40194 16730 40595
rect 17131 40470 20672 40595
rect 17131 40194 20670 40470
rect 16729 40193 17132 40194
rect 10849 17940 11411 17941
rect 10849 17380 10850 17940
rect 11410 17939 12672 17940
rect 11410 17381 12113 17939
rect 12671 17381 12672 17939
rect 11410 17380 12672 17381
rect 10849 17379 11411 17380
rect 25840 14539 26400 14540
rect 19064 14533 19624 14534
rect 12246 14461 12806 14462
rect 5522 14341 6082 14342
rect 5522 13783 5523 14341
rect 6081 13783 6082 14341
rect 5522 13702 6082 13783
rect 12246 13903 12247 14461
rect 12805 13903 12806 14461
rect 12246 13702 12806 13903
rect 19064 13975 19065 14533
rect 19623 13975 19624 14533
rect 19064 13820 19624 13975
rect 25840 13981 25841 14539
rect 26399 13981 26400 14539
rect 19064 13702 19650 13820
rect 4268 13142 7336 13702
rect 11016 13142 14084 13702
rect 17838 13142 20906 13702
rect 25840 13698 26400 13981
rect 24576 13138 27644 13698
rect 800 4035 1858 4036
rect 800 3637 1459 4035
rect 1857 3637 1858 4035
rect 800 3636 1858 3637
rect 800 1000 1200 3636
rect 19551 766 30599 767
rect 19551 486 19552 766
rect 19832 486 30599 766
rect 19551 485 30599 486
rect 30317 317 30599 485
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30358 114 30558 317
rect 30362 0 30542 114
use adc_digital_control  adc_digital_control_0
timestamp 1727826562
transform -1 0 22030 0 1 40330
box 514 0 4576 3000
use opamp_ladder  opamp_ladder_0
timestamp 1727841813
transform 0 -1 14726 1 0 -2498
box 3748 -14788 16764 11394
<< labels >>
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
