magic
tech sky130A
timestamp 1730259253
<< metal2 >>
rect 9600 1660 10140 1680
rect 9380 1640 10360 1660
rect 40 1540 560 1640
rect 4300 1620 4440 1640
rect 9240 1620 10480 1640
rect 4280 1600 4460 1620
rect 6300 1600 6560 1620
rect 9140 1600 10580 1620
rect 4260 1580 4480 1600
rect 6320 1580 6580 1600
rect 9120 1580 10660 1600
rect 4240 1560 4500 1580
rect 6300 1560 6600 1580
rect 9100 1560 10740 1580
rect 4220 1540 4520 1560
rect 40 960 580 1540
rect 4200 1520 4520 1540
rect 6300 1540 6620 1560
rect 9080 1540 10800 1560
rect 4200 1500 4540 1520
rect 6300 1500 6640 1540
rect 9060 1520 10860 1540
rect 9020 1500 10920 1520
rect 4180 1480 4560 1500
rect 6300 1480 6660 1500
rect 8960 1480 10960 1500
rect 4160 1460 4580 1480
rect 6300 1460 6680 1480
rect 8880 1460 11020 1480
rect 4140 1440 4600 1460
rect 6300 1440 6700 1460
rect 8840 1440 11060 1460
rect 1860 1420 2040 1440
rect 4120 1420 4620 1440
rect 6300 1420 6720 1440
rect 8780 1420 11100 1440
rect 1860 1400 2120 1420
rect 4100 1400 4640 1420
rect 6300 1400 6740 1420
rect 8740 1400 11140 1420
rect 1860 1380 2180 1400
rect 4080 1380 4660 1400
rect 6300 1380 6760 1400
rect 8700 1380 9640 1400
rect 9980 1380 11180 1400
rect 1860 1360 2220 1380
rect 4060 1360 4680 1380
rect 6300 1360 6780 1380
rect 8660 1360 9400 1380
rect 10200 1360 11200 1380
rect 1860 1340 2240 1360
rect 4040 1340 4700 1360
rect 6300 1340 6800 1360
rect 8620 1340 9260 1360
rect 10320 1340 11240 1360
rect 1860 1320 2280 1340
rect 4020 1320 4720 1340
rect 6300 1320 6820 1340
rect 8580 1320 9160 1340
rect 10420 1320 11280 1340
rect 1860 1300 2300 1320
rect 1860 1280 2320 1300
rect 4000 1280 4740 1320
rect 6300 1280 6840 1320
rect 8560 1300 9080 1320
rect 10500 1300 11300 1320
rect 8520 1280 9000 1300
rect 10560 1280 11320 1300
rect 1860 1260 2340 1280
rect 3980 1260 4760 1280
rect 6300 1260 6860 1280
rect 8500 1260 8940 1280
rect 10620 1260 11360 1280
rect 1860 1220 2360 1260
rect 3960 1240 4780 1260
rect 3940 1220 4800 1240
rect 1860 1200 2380 1220
rect 3920 1200 4172 1220
rect 4200 1200 4820 1220
rect 1860 1140 2400 1200
rect 3900 1180 4160 1200
rect 4220 1180 4840 1200
rect 3880 1160 4140 1180
rect 4240 1160 4860 1180
rect 3860 1140 4120 1160
rect 4260 1140 4880 1160
rect 40 940 600 960
rect 1860 940 2420 1140
rect 4280 1120 4900 1140
rect 4300 1100 4920 1120
rect 4320 1080 4940 1100
rect 4340 1060 4960 1080
rect 4360 1040 4960 1060
rect 4380 1020 4980 1040
rect 4400 1000 5000 1020
rect 4420 980 5020 1000
rect 4440 960 5040 980
rect 4460 940 5060 960
rect 40 920 720 940
rect 1840 920 2420 940
rect 4480 920 5080 940
rect 40 720 2420 920
rect 3640 912 4432 920
rect 3640 900 4452 912
rect 4480 900 5100 920
rect 3620 880 5120 900
rect 3600 860 5140 880
rect 3580 840 5160 860
rect 3560 820 5180 840
rect 3540 800 5180 820
rect 3520 780 5200 800
rect 3500 760 5220 780
rect 3480 740 5240 760
rect 40 700 740 720
rect 1840 700 2420 720
rect 3460 720 5260 740
rect 3460 700 5280 720
rect 60 100 740 700
rect 1860 100 2420 700
rect 3440 680 4040 700
rect 4680 680 5300 700
rect 3420 660 4020 680
rect 4700 660 5320 680
rect 3400 640 4000 660
rect 4720 640 5340 660
rect 3380 620 3980 640
rect 4740 620 5360 640
rect 3360 600 3960 620
rect 4760 600 5380 620
rect 3340 580 3940 600
rect 4780 580 5400 600
rect 3320 560 3920 580
rect 4800 560 5400 580
rect 3300 540 3900 560
rect 4820 540 5420 560
rect 3280 520 3880 540
rect 4820 520 5440 540
rect 3260 500 3860 520
rect 4840 500 5460 520
rect 3260 480 3840 500
rect 4860 480 5480 500
rect 6300 480 6880 1260
rect 8480 1240 8900 1260
rect 10680 1240 11380 1260
rect 8440 1220 8840 1240
rect 10720 1220 11400 1240
rect 8420 1200 8800 1220
rect 10760 1200 11420 1220
rect 8400 1180 8760 1200
rect 10780 1180 11440 1200
rect 8380 1160 8720 1180
rect 10820 1160 11460 1180
rect 8360 1140 8680 1160
rect 10860 1140 11480 1160
rect 8360 1120 8660 1140
rect 10880 1120 11480 1140
rect 8340 1100 8620 1120
rect 10900 1100 11500 1120
rect 8320 1080 8600 1100
rect 10920 1080 11520 1100
rect 8320 1060 8580 1080
rect 10940 1060 11520 1080
rect 8340 1040 8560 1060
rect 10960 1040 11540 1060
rect 8360 1020 8540 1040
rect 10980 1020 11540 1040
rect 8400 1000 8520 1020
rect 11000 1000 11560 1020
rect 8420 980 8500 1000
rect 8440 960 8500 980
rect 9680 960 9920 980
rect 11020 960 11580 1000
rect 9620 940 9980 960
rect 9580 920 10020 940
rect 11040 920 11600 960
rect 9540 900 10060 920
rect 11040 900 11660 920
rect 9520 880 10080 900
rect 9500 760 10100 880
rect 11060 780 11920 900
rect 11040 760 11920 780
rect 9520 740 10080 760
rect 11040 740 11900 760
rect 9540 720 10060 740
rect 11020 720 11600 740
rect 9560 700 10040 720
rect 11020 700 11580 720
rect 9600 680 10000 700
rect 11000 680 11580 700
rect 9640 660 9960 680
rect 11000 660 11560 680
rect 9740 640 9860 660
rect 10980 640 11560 660
rect 10960 620 11540 640
rect 10940 600 11520 620
rect 10920 580 11500 600
rect 10880 560 11500 580
rect 10860 540 11480 560
rect 10820 520 11460 540
rect 10800 500 11440 520
rect 10760 480 11420 500
rect 3240 460 3840 480
rect 4880 460 5500 480
rect 3220 440 3820 460
rect 4900 440 5520 460
rect 6300 440 6900 480
rect 10720 460 11400 480
rect 10680 440 11380 460
rect 3200 420 3800 440
rect 4920 420 5540 440
rect 6300 420 6920 440
rect 10640 420 11360 440
rect 3180 400 3780 420
rect 4940 400 5560 420
rect 6300 400 6940 420
rect 10580 400 11340 420
rect 3160 380 3760 400
rect 4960 380 5580 400
rect 6300 380 6980 400
rect 10520 380 11320 400
rect 3140 360 3740 380
rect 4980 360 5600 380
rect 6300 360 7040 380
rect 10460 360 11280 380
rect 3120 340 3720 360
rect 5000 340 5620 360
rect 3100 320 3700 340
rect 5020 320 5620 340
rect 6300 340 8180 360
rect 9040 340 9120 360
rect 10380 340 11260 360
rect 6300 320 8220 340
rect 9040 320 9240 340
rect 10280 320 11240 340
rect 3080 300 3680 320
rect 5040 300 5640 320
rect 6320 300 8240 320
rect 9040 300 9380 320
rect 10180 300 11200 320
rect 3060 280 3660 300
rect 5060 280 5660 300
rect 6320 280 8260 300
rect 9040 280 9580 300
rect 10040 280 11160 300
rect 3060 260 3640 280
rect 5080 260 5680 280
rect 6340 260 8300 280
rect 9040 260 11140 280
rect 3040 240 3620 260
rect 5080 240 5700 260
rect 6360 240 8320 260
rect 9040 240 11100 260
rect 3020 220 3600 240
rect 5100 220 5720 240
rect 6380 220 8340 240
rect 9040 220 11060 240
rect 3000 200 3580 220
rect 5120 200 5740 220
rect 6400 200 8380 220
rect 2980 180 3580 200
rect 5140 180 5760 200
rect 6420 180 8380 200
rect 9040 200 11020 220
rect 9040 180 10960 200
rect 2960 160 3560 180
rect 5160 160 5780 180
rect 6440 160 8380 180
rect 9080 160 10920 180
rect 2940 140 3540 160
rect 5180 140 5800 160
rect 6460 140 8380 160
rect 9180 140 10860 160
rect 2920 120 3520 140
rect 5200 120 5820 140
rect 6480 120 8380 140
rect 9320 120 10780 140
rect 5220 100 5300 120
rect 6500 100 7840 120
rect 9460 100 10700 120
rect 9560 80 10620 100
rect 9580 60 10520 80
rect 9600 40 10380 60
rect 9640 20 10180 40
<< end >>
