magic
tech sky130A
magscale 1 2
timestamp 1728774904
<< metal1 >>
rect 8796 3414 8862 3470
rect 8796 2676 8862 2732
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 8796 -656 8862 -600
rect 0 -1200 200 -1000
rect 8796 -1076 8862 -1020
rect 0 -1600 200 -1400
use sky130_fd_pr__pfet_01v8_XPP7BA  XM1
timestamp 1728771870
transform 1 0 7974 0 1 1241
box -256 -819 256 819
use sky130_fd_pr__pfet_01v8_XPP7BA  XM2
timestamp 1728771870
transform 1 0 8380 0 1 1241
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_3BHWKV  XM3
timestamp 1728771870
transform 1 0 7974 0 1 -388
box -256 -810 256 810
use sky130_fd_pr__nfet_01v8_3BHWKV  XM4
timestamp 1728771870
transform 1 0 8380 0 1 -388
box -256 -810 256 810
use sky130_fd_pr__pfet_01v8_XPP7BA  XM5
timestamp 1728771870
transform 1 0 8380 0 1 2773
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_848SAM  XM6
timestamp 1728771870
transform 1 0 8829 0 1 -838
box -211 -360 211 360
use sky130_fd_pr__pfet_01v8_XGSNAL  XM7
timestamp 1728771870
transform 1 0 8829 0 1 3073
box -211 -519 211 519
use sky130_fd_pr__pfet_01v8_XPP7BA  XM8
timestamp 1728771870
transform 1 0 7974 0 1 2773
box -256 -819 256 819
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR1
timestamp 1728771870
transform 0 -1 6736 1 0 -701
box -201 -982 201 982
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR2
timestamp 1728771870
transform 0 -1 6736 1 0 -405
box -201 -982 201 982
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR3
timestamp 1728771870
transform 0 -1 6736 1 0 -109
box -201 -982 201 982
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR4
timestamp 1728771870
transform 0 -1 6736 1 0 187
box -201 -982 201 982
use sky130_fd_pr__res_high_po_0p35_WFRDHL  XR
timestamp 1728771870
transform 0 -1 6736 1 0 -997
box -201 -982 201 982
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 vin_n
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 vin_p
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vout
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VGND
port 4 nsew
<< end >>
