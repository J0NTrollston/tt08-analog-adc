* Simulation of an R2R DAC with Verilator and d_cosim

.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* https://sourceforge.net/p/ngspice/ngspice/ci/master/tree/examples/xspice/verilator/

* The digital portion of the circuit is specified in compiled Verilog.
* list the inputs and outputs
adut [clk reset_n btn analog_to_digital_in_3 analog_to_digital_in_2 analog_to_digital_in_1 analog_to_digital_in_0 ] [encoded_out_1 encoded_out_0 control_2 control_1 control_0] null dut
.model dut d_cosim simulation="./adc_digital_control.so"

* connect the driver to the R2R dac
* had to edit spice exported by xschem to add the subckt and ends

.include "../xschem/simulation/opamp_ladder.spice" 
*.include "../mag/r2r.spice" 

xopamp_ladder vcc in0 0 analog_to_digital_in_3 analog_to_digital_in_2 analog_to_digital_in_1 analog_to_digital_in_0 opamp_ladder

* simulate tt output path
R1 out pin_out 500
C1 out 0 5p



**** End of the ADC and its subcircuits.  Begin test circuit ****

.param vcc=1.8
vcc vcc 0 {vcc}

* Digital clock signal

* aclock 0 clk clock
* .model clock d_osc cntl_array=[-1 1] freq_array=[1Meg 1Meg]

* reset signal
* Vreset n_rst 0 PULSE 3 0 1n 1u 10p 1u 500u

Vin0 in0 0 PULSE 0 1.8 50u 350u 1n



.control
 tran 100n 500u UIC
plot in0 analog_to_digital_in_0 analog_to_digital_in_1 analog_to_digital_in_2 analog_to_digital_in_3
plot in0 encoded_out_0 encoded_out_1
.endc
.end
