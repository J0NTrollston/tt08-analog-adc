magic
tech sky130A
magscale 1 2
timestamp 1727817497
<< error_s >>
rect 7274 8232 7280 8238
rect 7468 8232 7474 8238
rect 7268 8226 7274 8232
rect 7474 8226 7480 8232
rect 7268 8032 7274 8038
rect 7474 8032 7480 8038
rect 7274 8026 7280 8032
rect 7468 8026 7474 8032
rect 7270 1480 7276 1486
rect 7464 1480 7470 1486
rect 7264 1474 7270 1480
rect 7470 1474 7476 1480
rect 7264 1280 7270 1286
rect 7470 1280 7476 1286
rect 7270 1274 7276 1280
rect 7464 1274 7470 1280
rect 4108 -2566 4114 -2560
rect 4302 -2566 4308 -2560
rect 4102 -2572 4108 -2566
rect 4308 -2572 4314 -2566
rect 4102 -2766 4108 -2760
rect 4308 -2766 4314 -2760
rect 4108 -2772 4114 -2766
rect 4302 -2772 4308 -2766
rect 7274 -8910 7280 -8904
rect 7468 -8910 7474 -8904
rect 7268 -8916 7274 -8910
rect 7474 -8916 7480 -8910
rect 7268 -9110 7274 -9104
rect 7474 -9110 7480 -9104
rect 7274 -9116 7280 -9110
rect 7468 -9116 7474 -9110
<< pwell >>
rect 4630 11194 4806 11354
<< viali >>
rect 4906 8700 4940 10622
rect 4914 5932 4948 7854
rect 4940 -828 4974 1094
rect 4946 -7634 4980 -5712
rect 4954 -14380 4988 -12458
<< metal1 >>
rect 3830 11194 7690 11394
rect 4630 10518 4806 11194
rect 4894 10622 5087 10630
rect 4630 8386 4814 8804
rect 4894 8700 4906 10622
rect 4940 9774 5087 10622
rect 4940 9769 5188 9774
rect 4940 9768 5189 9769
rect 4940 9589 5009 9768
rect 5188 9589 5189 9768
rect 4940 9588 5189 9589
rect 4940 9583 5188 9588
rect 4940 8700 5087 9583
rect 4894 8692 5087 8700
rect 4630 8380 4832 8386
rect 4630 8180 4632 8380
rect 4630 8174 4832 8180
rect 4630 7750 4814 8174
rect 4902 7854 5094 7862
rect 4638 3660 4840 6036
rect 4902 5932 4914 7854
rect 4948 6983 5094 7854
rect 4948 6978 5195 6983
rect 4948 6977 5196 6978
rect 4948 6799 5017 6977
rect 5195 6799 5196 6977
rect 4948 6798 5196 6799
rect 4948 6793 5195 6798
rect 4948 5932 5094 6793
rect 4902 5924 5094 5932
rect 4632 3654 4840 3660
rect 4832 3454 4840 3654
rect 4632 3448 4840 3454
rect 4638 990 4840 3448
rect 5282 4642 5511 11194
rect 5834 9792 6062 9798
rect 5834 7002 6062 9564
rect 6600 8974 7470 9028
rect 6600 8846 7590 8974
rect 6600 8828 7470 8846
rect 5828 6774 5834 7002
rect 6062 6774 6068 7002
rect 5834 5716 6062 6774
rect 5828 5516 5834 5716
rect 6034 5516 6062 5716
rect 5482 4442 5511 4642
rect 4928 1094 5109 1102
rect 3748 -2766 4108 -2566
rect 4664 -3198 4846 -724
rect 4928 -828 4940 1094
rect 4974 215 5109 1094
rect 4974 209 5205 215
rect 4974 40 5036 209
rect 4974 34 5205 40
rect 4974 -828 5109 34
rect 4928 -836 5109 -828
rect 5282 -2182 5511 4442
rect 5834 238 6062 5516
rect 6600 2276 6828 8828
rect 7270 5716 7470 7426
rect 16350 6338 16736 6538
rect 7266 5516 7272 5716
rect 7472 5682 7478 5716
rect 7472 5518 7654 5682
rect 7472 5516 7478 5518
rect 7256 4442 7262 4642
rect 7462 4442 7468 4642
rect 6600 2076 7466 2276
rect 5828 10 5834 238
rect 6062 10 6068 238
rect 5834 -1036 6062 10
rect 5830 -1236 5836 -1036
rect 6036 -1236 6062 -1036
rect 5482 -2382 5511 -2182
rect 4664 -3204 4868 -3198
rect 4664 -3404 4668 -3204
rect 4664 -3410 4868 -3404
rect 4664 -5816 4846 -3410
rect 4934 -5712 5107 -5704
rect 4670 -9968 4854 -7530
rect 4934 -7634 4946 -5712
rect 4980 -6587 5107 -5712
rect 4980 -6593 5213 -6587
rect 4980 -6754 5052 -6593
rect 4980 -6760 5213 -6754
rect 4980 -7634 5107 -6760
rect 4934 -7642 5107 -7634
rect 5282 -8910 5511 -2382
rect 5834 -6560 6062 -1236
rect 6600 -4548 6828 2076
rect 7266 -1036 7466 674
rect 16350 -414 16728 -214
rect 7262 -1236 7268 -1036
rect 7468 -1236 7474 -1036
rect 7264 -2382 7270 -2182
rect 7470 -2382 7476 -2182
rect 6600 -4748 7474 -4548
rect 5828 -6788 5834 -6560
rect 6062 -6788 6068 -6560
rect 5834 -7860 6062 -6788
rect 5834 -8060 5838 -7860
rect 6038 -8060 6062 -7860
rect 5482 -9110 5512 -8910
rect 5282 -9116 5482 -9110
rect 4670 -9974 4870 -9968
rect 4670 -10174 4671 -9974
rect 4670 -10180 4870 -10174
rect 4670 -12562 4854 -10180
rect 4942 -12458 5127 -12450
rect 4678 -14586 4854 -14276
rect 4942 -14380 4954 -12458
rect 4988 -13344 5127 -12458
rect 5834 -13324 6062 -8060
rect 6600 -11276 6828 -4748
rect 7272 -5544 7278 -5344
rect 7478 -5544 7484 -5344
rect 7274 -7860 7474 -6150
rect 16348 -7238 16744 -7038
rect 7270 -8060 7276 -7860
rect 7476 -8060 7482 -7860
rect 7474 -9110 7642 -8910
rect 6600 -11330 7478 -11276
rect 6600 -11458 7606 -11330
rect 6600 -11476 7478 -11458
rect 6608 -12272 6614 -12072
rect 6814 -12272 7482 -12072
rect 4988 -13350 5220 -13344
rect 4988 -13525 5045 -13350
rect 4988 -13531 5220 -13525
rect 4988 -14380 5127 -13531
rect 5828 -13552 5834 -13324
rect 6062 -13552 6068 -13324
rect 4942 -14388 5127 -14380
rect 3792 -14622 4854 -14586
rect 5834 -14622 6062 -13552
rect 7278 -14622 7478 -12878
rect 16352 -13966 16764 -13766
rect 3792 -14786 7748 -14622
<< via1 >>
rect 5009 9589 5188 9768
rect 4632 8180 4832 8380
rect 5017 6799 5195 6977
rect 4632 3454 4832 3654
rect 5834 9564 6062 9792
rect 5834 6774 6062 7002
rect 5834 5516 6034 5716
rect 5282 4442 5482 4642
rect 4108 -2766 4308 -2566
rect 5036 40 5205 209
rect 7274 8032 7474 8232
rect 7272 5516 7472 5716
rect 7262 4442 7462 4642
rect 5834 10 6062 238
rect 5836 -1236 6036 -1036
rect 5282 -2382 5482 -2182
rect 4668 -3404 4868 -3204
rect 5052 -6754 5213 -6593
rect 7270 1280 7470 1480
rect 7268 -1236 7468 -1036
rect 7270 -2382 7470 -2182
rect 5834 -6788 6062 -6560
rect 5838 -8060 6038 -7860
rect 5282 -9110 5482 -8910
rect 4671 -10174 4870 -9974
rect 7278 -5544 7478 -5344
rect 7276 -8060 7476 -7860
rect 7274 -9110 7474 -8910
rect 6614 -12272 6814 -12072
rect 5045 -13525 5220 -13350
rect 5834 -13552 6062 -13324
<< metal2 >>
rect 5828 9768 5834 9792
rect 5003 9589 5009 9768
rect 5188 9589 5834 9768
rect 5828 9564 5834 9589
rect 6062 9564 6068 9792
rect 4626 8180 4632 8380
rect 4832 8232 6442 8380
rect 4832 8180 7274 8232
rect 6242 8032 7274 8180
rect 5834 7002 6062 7008
rect 5011 6799 5017 6977
rect 5195 6799 5834 6977
rect 5834 6768 6062 6774
rect 5834 5716 6034 5722
rect 7272 5716 7472 5722
rect 6034 5516 7272 5716
rect 5834 5510 6034 5516
rect 7272 5510 7472 5516
rect 7262 4642 7462 4648
rect 5276 4442 5282 4642
rect 5482 4442 7262 4642
rect 7262 4436 7462 4442
rect 4626 3454 4632 3654
rect 4832 3454 6442 3654
rect 6242 1480 6442 3454
rect 6242 1280 7270 1480
rect 5834 238 6062 244
rect 5030 40 5036 209
rect 5205 40 5834 209
rect 5834 4 6062 10
rect 5836 -1036 6036 -1030
rect 7268 -1036 7468 -1030
rect 6036 -1236 7268 -1036
rect 5836 -1242 6036 -1236
rect 7268 -1242 7468 -1236
rect 7270 -2182 7470 -2176
rect 5276 -2382 5282 -2182
rect 5482 -2382 7270 -2182
rect 7270 -2388 7470 -2382
rect 4308 -2766 6810 -2566
rect 4662 -3404 4668 -3204
rect 4868 -3404 6438 -3204
rect 6238 -5344 6438 -3404
rect 7278 -5344 7478 -5338
rect 6238 -5544 7278 -5344
rect 7278 -5550 7478 -5544
rect 5834 -6560 6062 -6554
rect 5046 -6754 5052 -6593
rect 5213 -6754 5834 -6593
rect 5834 -6794 6062 -6788
rect 7276 -7860 7476 -7854
rect 5832 -8060 5838 -7860
rect 6038 -8060 7276 -7860
rect 7276 -8066 7476 -8060
rect 5276 -9110 5282 -8910
rect 5482 -9110 7274 -8910
rect 4665 -10174 4671 -9974
rect 4870 -10174 6440 -9974
rect 6240 -12072 6440 -10174
rect 6614 -12072 6814 -12066
rect 6240 -12272 6614 -12072
rect 6614 -12278 6814 -12272
rect 5834 -13324 6062 -13318
rect 5039 -13525 5045 -13350
rect 5220 -13525 5834 -13350
rect 5834 -13558 6062 -13552
use opamp  x1
timestamp 1727813218
transform 1 0 4536 0 1 -12486
box 2738 -2302 11916 3576
use opamp  x2
timestamp 1727813218
transform 1 0 4532 0 1 -5758
box 2738 -2302 11916 3576
use opamp  x3
timestamp 1727813218
transform 1 0 4524 0 1 1066
box 2738 -2302 11916 3576
use opamp  x4
timestamp 1727813218
transform 1 0 4528 0 1 7818
box 2738 -2302 11916 3576
use sky130_fd_pr__res_generic_nd_BRW5P9  XR1
timestamp 1727813169
transform 1 0 4718 0 1 9661
box -258 -1101 258 1101
use sky130_fd_pr__res_generic_nd_BRW5P9  XR2
timestamp 1727813169
transform 1 0 4766 0 1 -13419
box -258 -1101 258 1101
use sky130_fd_pr__res_generic_nd_BRW5P9  XR3
timestamp 1727813169
transform 1 0 4758 0 1 -6673
box -258 -1101 258 1101
use sky130_fd_pr__res_generic_nd_BRW5P9  XR4
timestamp 1727813169
transform 1 0 4752 0 1 133
box -258 -1101 258 1101
use sky130_fd_pr__res_generic_nd_BRW5P9  XR5
timestamp 1727813169
transform 1 0 4726 0 1 6893
box -258 -1101 258 1101
<< labels >>
flabel metal1 3830 11194 4030 11394 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 3792 -14786 3992 -14586 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 3748 -2766 3948 -2566 0 FreeSans 256 0 0 0 in
port 1 nsew
flabel metal1 16564 -13966 16764 -13766 0 FreeSans 256 0 0 0 out0
port 6 nsew
flabel metal1 16544 -7238 16744 -7038 0 FreeSans 256 0 0 0 out1
port 5 nsew
flabel metal1 16528 -414 16728 -214 0 FreeSans 256 0 0 0 out2
port 4 nsew
flabel metal1 16536 6338 16736 6538 0 FreeSans 256 0 0 0 out3
port 3 nsew
<< end >>
