magic
tech sky130A
magscale 1 2
timestamp 1727469472
<< checkpaint >>
rect 9438 -103 12474 -50
rect 2290 -217 5322 -164
rect 2290 -4304 5781 -217
rect 9438 -482 12937 -103
rect 2749 -4357 5781 -4304
rect 8926 -4145 12937 -482
rect 8926 -4622 12884 -4145
rect 9385 -4675 12884 -4622
rect 9848 -4728 12884 -4675
<< error_p >>
rect 5392 1304 5962 1340
rect 4924 1242 5962 1304
rect 4924 1136 5004 1242
rect 5092 1172 5794 1242
rect 5092 1170 5674 1172
rect 5794 1170 5814 1172
rect 5932 1170 5962 1242
rect 5092 1052 5638 1170
rect 5202 1031 5638 1052
rect 4972 222 5004 390
<< error_s >>
rect 5202 1028 5638 1031
rect 5202 1024 5384 1028
rect 5506 1024 5638 1028
rect 5456 1004 5638 1024
rect 5336 222 5404 390
rect 5456 386 5590 1004
rect 5140 218 5172 222
rect 5236 218 5404 222
rect 5436 218 5590 386
rect 5236 -156 5322 -10
rect 5322 -178 5404 -156
rect 5456 -178 5576 98
rect 5604 -178 5624 218
rect 9416 -620 9616 -600
rect 10155 -620 10219 -257
rect 9436 -779 9437 -620
rect 9596 -779 9616 -620
rect 9436 -780 9616 -779
rect 10048 -780 10219 -620
rect 3073 -1370 3108 -1336
rect 3074 -1389 3108 -1370
rect 2926 -2136 2944 -2102
rect 2954 -2136 2972 -2074
rect 2926 -2302 2944 -2300
rect 2954 -2330 2972 -2300
rect 3093 -2902 3108 -1389
rect 3127 -1423 3162 -1389
rect 3532 -1423 3567 -1406
rect 3127 -2902 3161 -1423
rect 3533 -1424 3567 -1423
rect 3533 -1460 3603 -1424
rect 3550 -1494 3621 -1460
rect 3991 -1494 4026 -1460
rect 3127 -2936 3142 -2902
rect 3550 -2955 3620 -1494
rect 3992 -1513 4026 -1494
rect 4468 -1513 4521 -1512
rect 3844 -2136 3858 -1772
rect 3872 -2136 3886 -1744
rect 3550 -2991 3603 -2955
rect 4011 -3008 4026 -1513
rect 4045 -1547 4080 -1513
rect 4450 -1547 4521 -1513
rect 4045 -3008 4079 -1547
rect 4451 -1548 4521 -1547
rect 4468 -1582 4539 -1548
rect 4900 -1565 4980 -1512
rect 4045 -3042 4060 -3008
rect 4468 -3061 4538 -1582
rect 4900 -1766 5092 -1565
rect 5368 -1635 5403 -1601
rect 5369 -1654 5403 -1635
rect 4900 -1784 5099 -1766
rect 4900 -1794 5092 -1784
rect 4762 -2136 4776 -1794
rect 4790 -2136 4804 -1794
rect 4468 -3097 4521 -3061
rect 4929 -3114 4944 -1794
rect 4963 -3114 4997 -1794
rect 5077 -1834 5111 -1796
rect 5236 -1806 5384 -1762
rect 5255 -1834 5289 -1806
rect 5388 -1834 5403 -1654
rect 5422 -1688 5457 -1654
rect 5422 -1834 5456 -1688
rect 5077 -1849 5736 -1834
rect 5077 -1894 5748 -1849
rect 5077 -1946 5111 -1894
rect 5255 -1946 5289 -1894
rect 5048 -1980 5289 -1946
rect 5077 -2972 5111 -1980
rect 5255 -2972 5289 -1980
rect 4963 -3148 4978 -3114
rect 5388 -3167 5403 -1894
rect 5422 -3167 5456 -1894
rect 5536 -1934 5570 -1894
rect 5714 -1934 5748 -1894
rect 5536 -2050 5800 -1934
rect 5536 -3025 5570 -2050
rect 5714 -3025 5748 -2050
rect 5828 -2689 5862 -2671
rect 5828 -2725 5898 -2689
rect 5845 -2759 5916 -2725
rect 5422 -3201 5437 -3167
rect 5845 -3220 5915 -2759
rect 5845 -3256 5898 -3220
rect 10155 -3281 10219 -780
rect 11143 -1380 11178 -1346
rect 11144 -1399 11178 -1380
rect 11163 -2796 11178 -1399
rect 11197 -1433 11232 -1399
rect 11197 -2796 11231 -1433
rect 11197 -2830 11212 -2796
<< nwell >>
rect 5004 1172 5932 1242
rect 5004 1170 5560 1172
rect 5794 1170 5932 1172
rect 5004 1136 5932 1170
rect 5004 1052 5092 1136
rect 5238 1052 5932 1136
rect 5004 1028 5932 1052
rect 5004 1024 5336 1028
rect 5506 1024 5932 1028
rect 5004 1004 5384 1024
rect 5004 222 5336 1004
rect 5004 218 5140 222
rect 5236 218 5336 222
rect 5456 218 5932 1024
rect 5236 -178 5322 -156
rect 5456 -178 5604 218
<< pwell >>
rect 5104 -524 5288 -518
rect 5104 -576 5304 -524
rect 5288 -584 5304 -576
rect 5456 -604 5552 -514
rect 4932 -1102 5092 -618
rect 5336 -660 5338 -620
rect 5456 -678 5604 -604
rect 5456 -758 5552 -678
rect 4900 -1794 5092 -1102
rect 5236 -1806 5384 -1762
rect 7844 -1796 7998 -620
rect 5104 -1894 5736 -1834
rect 5552 -2050 5800 -1934
<< viali >>
rect 5070 3064 5258 3098
rect 3546 1636 3580 2994
rect 6718 1738 6752 2996
rect 5048 1172 5280 1206
rect 5560 1172 5792 1206
rect 3548 -354 3582 888
rect 3548 -1876 3582 -634
rect 6502 -672 6734 -638
rect 5048 -1980 5280 -1946
rect 5560 -1980 5792 -1946
rect 7656 -1982 7888 -1948
<< metal1 >>
rect 2738 3376 6770 3576
rect 3522 2994 3678 3376
rect 3522 1636 3546 2994
rect 3580 2904 3678 2994
rect 3738 3012 3794 3018
rect 3738 2950 3794 2956
rect 4548 2904 4748 3376
rect 5064 3098 5264 3376
rect 5064 3064 5070 3098
rect 5258 3064 5264 3098
rect 5064 3052 5264 3064
rect 5136 3006 5192 3012
rect 5136 2944 5192 2950
rect 6558 2996 6770 3376
rect 9048 3130 9466 3294
rect 9630 3130 9636 3294
rect 5441 2904 5607 2905
rect 3580 2725 3700 2904
rect 3580 1726 3694 2725
rect 3838 1854 3952 2904
rect 3832 1734 4250 1854
rect 3838 1728 3952 1734
rect 3580 1636 3678 1726
rect 3522 1332 3678 1636
rect 3706 1618 3740 1674
rect 3796 1618 3826 1674
rect 2742 1156 2942 1210
rect 3522 1176 3848 1332
rect 2742 1131 3206 1156
rect 2742 1053 3103 1131
rect 3181 1053 3206 1131
rect 3692 1064 3848 1176
rect 2742 1028 3206 1053
rect 2742 1010 2942 1028
rect 3682 948 3852 1064
rect 3330 888 3594 896
rect 2746 394 2946 414
rect 2746 377 3226 394
rect 2746 259 3091 377
rect 3209 259 3226 377
rect 2746 243 3226 259
rect 2746 214 2946 243
rect 3330 -354 3548 888
rect 3582 -354 3594 888
rect 3682 784 3858 948
rect 3682 778 3852 784
rect 2742 -416 2942 -392
rect 3060 -416 3236 -410
rect 2742 -592 3060 -416
rect 3060 -598 3236 -592
rect 3330 -634 3594 -354
rect 3330 -1876 3548 -634
rect 3582 -1876 3594 -634
rect 3682 -416 3858 -250
rect 4130 -442 4250 1734
rect 4548 1726 5092 2904
rect 5236 1726 5607 2904
rect 5136 1680 5192 1686
rect 5136 1618 5192 1624
rect 4462 1544 4468 1600
rect 4524 1544 4530 1600
rect 3858 -562 4250 -442
rect 3682 -738 3858 -592
rect 4468 -626 4524 1544
rect 5441 1457 5607 1726
rect 6558 1738 6718 2996
rect 6752 2906 6770 2996
rect 6914 3006 6970 3012
rect 6914 2944 6970 2950
rect 9048 2906 9212 3130
rect 6752 1738 6866 2906
rect 7004 2742 9212 2906
rect 7004 2350 7168 2742
rect 6558 1730 6866 1738
rect 4724 1291 6120 1457
rect 4725 1012 4891 1291
rect 5040 1206 5288 1291
rect 5040 1172 5048 1206
rect 5280 1172 5288 1206
rect 5040 1160 5288 1172
rect 5552 1206 5800 1291
rect 5552 1172 5560 1206
rect 5792 1172 5800 1206
rect 5552 1160 5800 1172
rect 5136 1120 5192 1126
rect 5104 1064 5136 1120
rect 5192 1064 5224 1120
rect 5616 1064 5648 1120
rect 5704 1064 5736 1120
rect 5136 1058 5192 1064
rect 4725 -166 5092 1012
rect 5230 1004 5384 1024
rect 5236 21 5384 1004
rect 5230 -166 5384 21
rect 4725 -167 4891 -166
rect 5236 -178 5384 -166
rect 5104 -274 5136 -218
rect 5192 -274 5224 -218
rect 5288 -518 5384 -178
rect 5104 -576 5135 -518
rect 5193 -576 5384 -518
rect 5288 -604 5384 -576
rect 4612 -626 5092 -618
rect 4468 -682 5092 -626
rect 3330 -1884 3594 -1876
rect 2744 -2136 2944 -2102
rect 3330 -2136 3582 -1884
rect 3682 -2136 3858 -1772
rect 4612 -1794 5092 -682
rect 5236 -1652 5384 -604
rect 4612 -2136 4776 -1794
rect 5230 -1834 5384 -1652
rect 5456 -178 5604 1024
rect 5953 1012 6119 1291
rect 5748 -166 6119 1012
rect 5953 -167 6119 -166
rect 5456 -324 5552 -178
rect 6558 -200 6679 1730
rect 7010 1728 7168 2350
rect 6914 1680 6970 1686
rect 6914 1618 6970 1624
rect 5648 -218 5704 -212
rect 6558 -260 6588 -200
rect 6648 -260 6679 -200
rect 6558 -266 6679 -260
rect 7008 -92 7184 -86
rect 5648 -280 5704 -274
rect 7008 -310 7184 -268
rect 6194 -324 6546 -310
rect 5456 -352 6546 -324
rect 5456 -453 6100 -352
rect 6201 -453 6546 -352
rect 5456 -471 6546 -453
rect 5456 -604 5552 -471
rect 6194 -486 6546 -471
rect 6690 -486 7184 -310
rect 5647 -518 5705 -512
rect 5647 -582 5705 -576
rect 6588 -532 6648 -526
rect 7712 -576 7744 -520
rect 7800 -576 7832 -520
rect 6588 -598 6648 -592
rect 5456 -606 5604 -604
rect 5456 -1794 5608 -606
rect 5748 -626 6244 -618
rect 5748 -638 6742 -626
rect 5748 -672 6502 -638
rect 6734 -672 6742 -638
rect 5748 -754 6742 -672
rect 5748 -1794 6244 -754
rect 5104 -1894 5736 -1834
rect 5040 -1946 5288 -1934
rect 5040 -1980 5048 -1946
rect 5280 -1980 5288 -1946
rect 5040 -2136 5288 -1980
rect 5552 -1946 5800 -1934
rect 5552 -1980 5560 -1946
rect 5792 -1980 5800 -1946
rect 5552 -2136 5800 -1980
rect 6080 -2136 6244 -1794
rect 7430 -1796 7700 -620
rect 7838 -780 8574 -620
rect 8734 -780 8740 -620
rect 7844 -1796 7998 -780
rect 11716 -1320 11916 -1280
rect 11088 -1480 11094 -1320
rect 11254 -1480 11916 -1320
rect 7430 -1936 7614 -1796
rect 7712 -1896 7744 -1840
rect 7800 -1896 7832 -1840
rect 7430 -1948 7896 -1936
rect 7430 -1982 7656 -1948
rect 7888 -1982 7896 -1948
rect 7430 -2136 7896 -1982
rect 2744 -2300 8148 -2136
rect 2744 -2302 2944 -2300
<< via1 >>
rect 3738 2956 3794 3012
rect 5136 2950 5192 3006
rect 9466 3130 9630 3294
rect 3740 1618 3796 1674
rect 3103 1053 3181 1131
rect 3091 259 3209 377
rect 3060 -592 3236 -416
rect 3682 -592 3858 -416
rect 5136 1624 5192 1680
rect 4468 1544 4524 1600
rect 6914 2950 6970 3006
rect 5136 1064 5192 1120
rect 5648 1064 5704 1120
rect 5136 -274 5192 -218
rect 5135 -576 5193 -518
rect 6914 1624 6970 1680
rect 5648 -274 5704 -218
rect 6588 -260 6648 -200
rect 7008 -268 7184 -92
rect 6100 -453 6201 -352
rect 5647 -576 5705 -518
rect 6588 -592 6648 -532
rect 7744 -576 7800 -520
rect 8574 -780 8734 -620
rect 11094 -1480 11254 -1320
rect 7744 -1896 7800 -1840
<< metal2 >>
rect 9466 3294 9630 3300
rect 9630 3130 10006 3294
rect 10170 3130 10179 3294
rect 9466 3124 9630 3130
rect 3732 2956 3738 3012
rect 3794 2956 4098 3012
rect 4042 2346 4098 2956
rect 4828 2950 5136 3006
rect 5192 2950 6914 3006
rect 6970 2950 6976 3006
rect 4828 2346 4884 2950
rect 4042 2290 4884 2346
rect 3740 1674 3796 1680
rect 4042 1674 4098 2290
rect 3796 1618 4098 1674
rect 3740 1612 3796 1618
rect 4468 1600 4524 2290
rect 4828 1680 4884 2290
rect 4828 1624 5136 1680
rect 5192 1624 6914 1680
rect 6970 1624 6976 1680
rect 4468 1538 4524 1544
rect 3103 1216 3181 1227
rect 3103 1160 5448 1216
rect 3103 1131 3181 1160
rect 3103 1047 3181 1053
rect 3248 1120 3328 1132
rect 5392 1120 5448 1160
rect 5648 1120 5704 1126
rect 3248 1064 5136 1120
rect 5192 1064 5198 1120
rect 5392 1064 5648 1120
rect 3248 377 3328 1064
rect 3085 259 3091 377
rect 3209 259 3346 377
rect 4880 -218 4936 1064
rect 5136 -218 5192 -212
rect 4880 -274 5136 -218
rect 5392 -218 5448 1064
rect 5648 1058 5704 1064
rect 7008 304 7184 313
rect 7008 -92 7184 128
rect 5392 -274 5648 -218
rect 5704 -274 5710 -218
rect 6582 -260 6588 -200
rect 6648 -260 6852 -200
rect 5136 -280 5192 -274
rect 6100 -352 6201 -346
rect 3054 -592 3060 -416
rect 3236 -592 3682 -416
rect 3858 -592 3864 -416
rect 5135 -518 5193 -512
rect 5193 -576 5647 -518
rect 5705 -576 5711 -518
rect 5135 -582 5193 -576
rect 6100 -833 6201 -453
rect 6792 -532 6852 -260
rect 7002 -268 7008 -92
rect 7184 -268 7190 -92
rect 7744 -520 7800 -514
rect 6582 -592 6588 -532
rect 6648 -592 6852 -532
rect 7352 -576 7744 -520
rect 6100 -934 6501 -833
rect 6412 -1186 6488 -934
rect 7352 -1186 7408 -576
rect 7744 -582 7800 -576
rect 8574 -620 8734 -614
rect 8734 -780 9436 -620
rect 9596 -780 9605 -620
rect 8574 -786 8734 -780
rect 11094 -1089 11254 -1084
rect 6412 -1262 7408 -1186
rect 11090 -1239 11099 -1089
rect 11249 -1239 11258 -1089
rect 7352 -1840 7408 -1262
rect 11094 -1320 11254 -1239
rect 11094 -1486 11254 -1480
rect 7744 -1840 7800 -1834
rect 7352 -1896 7744 -1840
rect 7744 -1902 7800 -1896
<< via2 >>
rect 10006 3130 10170 3294
rect 7008 128 7184 304
rect 9436 -780 9596 -620
rect 11099 -1239 11249 -1089
<< metal3 >>
rect 10001 3294 10175 3299
rect 10001 3130 10006 3294
rect 10170 3130 10490 3294
rect 10654 3130 10660 3294
rect 10001 3125 10175 3130
rect 7008 754 7184 760
rect 7008 309 7184 578
rect 7003 304 7189 309
rect 7003 128 7008 304
rect 7184 128 7189 304
rect 7003 123 7189 128
rect 9431 -620 9601 -615
rect 9431 -780 9436 -620
rect 9596 -780 10048 -620
rect 10208 -780 10214 -620
rect 9431 -785 9601 -780
rect 11094 -875 11254 -874
rect 11089 -1033 11095 -875
rect 11253 -1033 11259 -875
rect 11094 -1089 11254 -1033
rect 11094 -1239 11099 -1089
rect 11249 -1239 11254 -1089
rect 11094 -1244 11254 -1239
<< via3 >>
rect 10490 3130 10654 3294
rect 7008 578 7184 754
rect 10048 -780 10208 -620
rect 11095 -1033 11253 -875
<< metal4 >>
rect 10489 3294 10655 3295
rect 10489 3130 10490 3294
rect 10654 3130 11254 3294
rect 10489 3129 10655 3130
rect 11090 1968 11254 3130
rect 7007 754 7185 755
rect 7007 578 7008 754
rect 7184 578 8366 754
rect 7007 577 7185 578
rect 10047 -620 10209 -619
rect 11094 -620 11254 368
rect 10047 -780 10048 -620
rect 10208 -780 11254 -620
rect 10047 -781 10209 -780
rect 11094 -875 11254 -780
rect 11094 -1033 11095 -875
rect 11253 -1033 11254 -875
rect 11094 -1034 11254 -1033
use sky130_fd_pr__cap_mim_m3_1_X5Y7W8  XC1
timestamp 1727401017
transform 1 0 8298 0 1 -1769
box -1941 -1540 1941 1540
use sky130_fd_pr__pfet_01v8_XPP7BA  XM1
timestamp 1727401017
transform 1 0 2888 0 1 -2119
box -256 -819 256 819
use sky130_fd_pr__pfet_01v8_XPP7BA  XM2
timestamp 1727401017
transform 1 0 3347 0 1 -2172
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_3BHWKV  XM3
timestamp 1727401017
transform 1 0 3806 0 1 -2234
box -256 -810 256 810
use sky130_fd_pr__nfet_01v8_3BHWKV  XM4
timestamp 1727401017
transform 1 0 4265 0 1 -2287
box -256 -810 256 810
use sky130_fd_pr__pfet_01v8_XPP7BA  XM5
timestamp 1727401017
transform 1 0 4724 0 1 -2331
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_3BHWKV  XM6
timestamp 1727401017
transform 1 0 10442 0 1 -2552
box -256 -810 256 810
use sky130_fd_pr__pfet_01v8_XPP7BA  XM7
timestamp 1727401017
transform 1 0 5183 0 1 -2384
box -256 -819 256 819
use sky130_fd_pr__pfet_01v8_XPP7BA  XM8
timestamp 1727401017
transform 1 0 5642 0 1 -2437
box -256 -819 256 819
use sky130_fd_pr__nfet_01v8_7QHW3M  XM9
timestamp 1727401017
transform 1 0 6101 0 1 -2999
box -256 -310 256 310
use sky130_fd_pr__res_generic_nd_GV5DH4  XR1
timestamp 1727401017
transform 1 0 10903 0 1 -2654
box -258 -761 258 761
use sky130_fd_pr__res_generic_nd_GV5DH4  XR2
timestamp 1727401017
transform 1 0 11366 0 1 -2707
box -258 -761 258 761
<< labels >>
flabel metal1 2742 -592 2942 -392 0 FreeSans 256 0 0 0 ZREF
port 1 nsew
flabel metal1 2744 -2302 2944 -2102 0 FreeSans 256 0 0 0 VGND
port 5 nsew
flabel metal1 2742 1010 2942 1210 0 FreeSans 256 0 0 0 vin_p
port 3 nsew
flabel metal1 2746 214 2946 414 0 FreeSans 256 0 0 0 vin_n
port 2 nsew
flabel metal1 2738 3376 2938 3576 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 11716 -1480 11916 -1280 0 FreeSans 256 0 0 0 Vout
port 4 nsew
<< end >>
