magic
tech sky130A
timestamp 1728462029
<< metal2 >>
rect 55000 102000 62000 103000
rect 54000 101000 63000 102000
rect 54000 100000 64000 101000
rect 53000 99000 64000 100000
rect 53000 98000 65000 99000
rect 52000 97000 65000 98000
rect 51000 96000 66000 97000
rect 51000 95000 67000 96000
rect 50000 94000 67000 95000
rect 50000 93000 68000 94000
rect 49000 92000 68000 93000
rect 49000 91000 69000 92000
rect 48000 90000 69000 91000
rect 210000 90000 214000 91000
rect 47000 89000 70000 90000
rect 207000 89000 217000 90000
rect 47000 88000 71000 89000
rect 206000 88000 218000 89000
rect 46000 87000 71000 88000
rect 46000 86000 58000 87000
rect 59000 86000 72000 87000
rect 205000 86000 219000 88000
rect 45000 85000 58000 86000
rect 60000 85000 72000 86000
rect 45000 84000 57000 85000
rect 60000 84000 73000 85000
rect 44000 83000 56000 84000
rect 61000 83000 73000 84000
rect 43000 82000 56000 83000
rect 62000 82000 74000 83000
rect 43000 81000 55000 82000
rect 62000 81000 75000 82000
rect 42000 80000 55000 81000
rect 63000 80000 75000 81000
rect 42000 79000 54000 80000
rect 63000 79000 76000 80000
rect 41000 78000 53000 79000
rect 40000 77000 53000 78000
rect 64000 78000 76000 79000
rect 64000 77000 77000 78000
rect 40000 76000 52000 77000
rect 65000 76000 77000 77000
rect 39000 75000 52000 76000
rect 66000 75000 78000 76000
rect 39000 74000 51000 75000
rect 66000 74000 79000 75000
rect 38000 73000 51000 74000
rect 67000 73000 79000 74000
rect 38000 72000 50000 73000
rect 67000 72000 80000 73000
rect 37000 71000 49000 72000
rect 68000 71000 80000 72000
rect 36000 70000 49000 71000
rect 36000 69000 48000 70000
rect 35000 68000 48000 69000
rect 53000 68000 65000 71000
rect 69000 70000 81000 71000
rect 69000 69000 82000 70000
rect 70000 68000 82000 69000
rect 35000 67000 47000 68000
rect 53000 67000 64000 68000
rect 70000 67000 83000 68000
rect 34000 66000 47000 67000
rect 52000 66000 64000 67000
rect 71000 66000 83000 67000
rect 34000 65000 46000 66000
rect 33000 64000 45000 65000
rect 52000 64000 63000 66000
rect 71000 65000 84000 66000
rect 72000 64000 84000 65000
rect 32000 63000 45000 64000
rect 51000 63000 63000 64000
rect 73000 63000 85000 64000
rect 32000 62000 44000 63000
rect 31000 61000 44000 62000
rect 51000 61000 62000 63000
rect 73000 62000 86000 63000
rect 74000 61000 86000 62000
rect 31000 60000 43000 61000
rect 51000 60000 61000 61000
rect 74000 60000 87000 61000
rect 30000 59000 43000 60000
rect 30000 58000 42000 59000
rect 50000 58000 61000 60000
rect 75000 59000 87000 60000
rect 137000 59000 149000 84000
rect 169000 59000 181000 84000
rect 204000 80000 220000 86000
rect 205000 78000 219000 80000
rect 206000 77000 218000 78000
rect 207000 76000 217000 77000
rect 209000 75000 215000 76000
rect 256000 70000 270000 71000
rect 193000 61000 219000 70000
rect 253000 69000 287000 70000
rect 251000 68000 287000 69000
rect 250000 67000 287000 68000
rect 248000 66000 287000 67000
rect 247000 64000 287000 66000
rect 246000 63000 287000 64000
rect 245000 62000 287000 63000
rect 245000 61000 259000 62000
rect 267000 61000 287000 62000
rect 296000 66000 308000 89000
rect 394000 82000 408000 84000
rect 434000 82000 447000 84000
rect 394000 81000 409000 82000
rect 395000 78000 409000 81000
rect 433000 80000 447000 82000
rect 433000 78000 446000 80000
rect 507000 79000 533000 89000
rect 574000 84000 579000 85000
rect 571000 83000 579000 84000
rect 567000 82000 579000 83000
rect 396000 75000 410000 78000
rect 432000 77000 446000 78000
rect 432000 75000 445000 77000
rect 397000 71000 411000 75000
rect 431000 74000 445000 75000
rect 431000 71000 444000 74000
rect 315000 70000 327000 71000
rect 313000 69000 329000 70000
rect 311000 68000 331000 69000
rect 398000 68000 412000 71000
rect 310000 67000 332000 68000
rect 309000 66000 333000 67000
rect 296000 64000 334000 66000
rect 399000 65000 413000 68000
rect 430000 67000 443000 71000
rect 466000 70000 481000 71000
rect 463000 69000 484000 70000
rect 461000 68000 486000 69000
rect 459000 67000 488000 68000
rect 400000 64000 413000 65000
rect 429000 64000 442000 67000
rect 458000 66000 489000 67000
rect 457000 65000 490000 66000
rect 456000 64000 491000 65000
rect 296000 61000 335000 64000
rect 400000 62000 414000 64000
rect 75000 58000 88000 59000
rect 29000 57000 41000 58000
rect 50000 57000 60000 58000
rect 76000 57000 88000 58000
rect 28000 56000 41000 57000
rect 28000 55000 40000 56000
rect 27000 54000 40000 55000
rect 49000 55000 60000 57000
rect 77000 56000 89000 57000
rect 77000 55000 90000 56000
rect 27000 53000 39000 54000
rect 49000 53000 59000 55000
rect 78000 54000 90000 55000
rect 78000 53000 91000 54000
rect 26000 52000 38000 53000
rect 25000 51000 38000 52000
rect 25000 50000 37000 51000
rect 24000 49000 37000 50000
rect 48000 50000 58000 53000
rect 68000 52000 70000 53000
rect 66000 51000 70000 52000
rect 79000 52000 91000 53000
rect 79000 51000 92000 52000
rect 64000 50000 69000 51000
rect 80000 50000 92000 51000
rect 48000 49000 57000 50000
rect 62000 49000 69000 50000
rect 24000 48000 36000 49000
rect 23000 47000 36000 48000
rect 47000 47000 57000 49000
rect 60000 48000 69000 49000
rect 81000 49000 93000 50000
rect 137000 49000 181000 59000
rect 81000 48000 94000 49000
rect 58000 47000 68000 48000
rect 23000 46000 35000 47000
rect 47000 46000 68000 47000
rect 82000 47000 94000 48000
rect 82000 46000 95000 47000
rect 22000 45000 34000 46000
rect 21000 44000 34000 45000
rect 46000 44000 68000 46000
rect 83000 45000 95000 46000
rect 84000 44000 96000 45000
rect 21000 43000 33000 44000
rect 20000 42000 33000 43000
rect 46000 42000 67000 44000
rect 84000 43000 97000 44000
rect 20000 41000 32000 42000
rect 19000 40000 32000 41000
rect 45000 41000 58000 42000
rect 45000 40000 55000 41000
rect 59000 40000 67000 42000
rect 85000 42000 97000 43000
rect 85000 41000 98000 42000
rect 86000 40000 98000 41000
rect 19000 39000 31000 40000
rect 45000 39000 53000 40000
rect 59000 39000 66000 40000
rect 86000 39000 99000 40000
rect 18000 38000 30000 39000
rect 45000 38000 51000 39000
rect 17000 37000 30000 38000
rect 44000 37000 49000 38000
rect 58000 37000 66000 39000
rect 87000 38000 99000 39000
rect 88000 37000 100000 38000
rect 17000 36000 29000 37000
rect 44000 36000 47000 37000
rect 16000 35000 29000 36000
rect 16000 34000 28000 35000
rect 58000 34000 65000 37000
rect 88000 36000 101000 37000
rect 89000 35000 101000 36000
rect 89000 34000 102000 35000
rect 15000 33000 28000 34000
rect 57000 33000 65000 34000
rect 90000 33000 102000 34000
rect 15000 32000 27000 33000
rect 14000 31000 26000 32000
rect 13000 30000 26000 31000
rect 57000 30000 64000 33000
rect 90000 32000 103000 33000
rect 91000 31000 103000 32000
rect 92000 30000 104000 31000
rect 13000 29000 25000 30000
rect 12000 28000 25000 29000
rect 57000 28000 63000 30000
rect 92000 29000 105000 30000
rect 12000 27000 24000 28000
rect 52000 27000 54000 28000
rect 11000 26000 23000 27000
rect 52000 26000 55000 27000
rect 56000 26000 63000 28000
rect 93000 28000 105000 29000
rect 93000 27000 106000 28000
rect 94000 26000 106000 27000
rect 10000 25000 23000 26000
rect 10000 24000 22000 25000
rect 9000 23000 22000 24000
rect 53000 24000 62000 26000
rect 65000 25000 66000 26000
rect 94000 25000 107000 26000
rect 63000 24000 66000 25000
rect 95000 24000 107000 25000
rect 9000 22000 21000 23000
rect 53000 22000 65000 24000
rect 96000 23000 108000 24000
rect 96000 22000 109000 23000
rect 137000 22000 149000 49000
rect 169000 22000 181000 49000
rect 206000 32000 219000 61000
rect 244000 60000 258000 61000
rect 268000 60000 281000 61000
rect 244000 59000 257000 60000
rect 269000 59000 281000 60000
rect 296000 60000 318000 61000
rect 320000 60000 336000 61000
rect 296000 59000 315000 60000
rect 322000 59000 336000 60000
rect 244000 57000 256000 59000
rect 244000 52000 255000 57000
rect 270000 56000 282000 59000
rect 271000 53000 282000 56000
rect 244000 50000 256000 52000
rect 270000 50000 282000 53000
rect 244000 48000 257000 50000
rect 269000 49000 282000 50000
rect 296000 58000 314000 59000
rect 296000 57000 313000 58000
rect 323000 57000 336000 59000
rect 401000 60000 414000 62000
rect 428000 61000 441000 64000
rect 455000 63000 492000 64000
rect 454000 62000 492000 63000
rect 454000 61000 493000 62000
rect 428000 60000 440000 61000
rect 453000 60000 472000 61000
rect 474000 60000 493000 61000
rect 401000 58000 415000 60000
rect 296000 56000 312000 57000
rect 296000 55000 311000 56000
rect 296000 54000 310000 55000
rect 296000 53000 309000 54000
rect 268000 48000 281000 49000
rect 245000 47000 259000 48000
rect 267000 47000 281000 48000
rect 245000 46000 281000 47000
rect 246000 45000 280000 46000
rect 247000 44000 279000 45000
rect 247000 43000 278000 44000
rect 246000 42000 277000 43000
rect 245000 41000 276000 42000
rect 245000 40000 275000 41000
rect 244000 39000 273000 40000
rect 244000 38000 255000 39000
rect 257000 38000 269000 39000
rect 243000 34000 254000 38000
rect 243000 33000 256000 34000
rect 243000 32000 258000 33000
rect 191000 22000 233000 32000
rect 243000 31000 275000 32000
rect 243000 30000 278000 31000
rect 244000 29000 281000 30000
rect 244000 28000 282000 29000
rect 245000 27000 284000 28000
rect 246000 25000 285000 27000
rect 245000 24000 286000 25000
rect 244000 23000 286000 24000
rect 243000 22000 257000 23000
rect 267000 22000 287000 23000
rect 296000 22000 308000 53000
rect 324000 22000 336000 57000
rect 402000 57000 415000 58000
rect 427000 58000 440000 60000
rect 452000 59000 469000 60000
rect 478000 59000 494000 60000
rect 452000 58000 467000 59000
rect 479000 58000 494000 59000
rect 427000 57000 439000 58000
rect 452000 57000 466000 58000
rect 480000 57000 495000 58000
rect 402000 55000 416000 57000
rect 403000 53000 416000 55000
rect 426000 54000 439000 57000
rect 451000 55000 465000 57000
rect 481000 56000 495000 57000
rect 482000 55000 495000 56000
rect 451000 54000 464000 55000
rect 426000 53000 438000 54000
rect 403000 52000 417000 53000
rect 404000 50000 417000 52000
rect 425000 51000 438000 53000
rect 450000 53000 464000 54000
rect 482000 53000 496000 55000
rect 425000 50000 437000 51000
rect 404000 48000 418000 50000
rect 405000 46000 418000 48000
rect 424000 48000 437000 50000
rect 424000 46000 436000 48000
rect 405000 45000 419000 46000
rect 406000 42000 419000 45000
rect 423000 45000 436000 46000
rect 450000 47000 463000 53000
rect 450000 45000 462000 47000
rect 423000 43000 435000 45000
rect 407000 39000 420000 42000
rect 422000 41000 435000 43000
rect 422000 39000 434000 41000
rect 408000 38000 434000 39000
rect 450000 39000 463000 45000
rect 483000 40000 496000 53000
rect 482000 39000 496000 40000
rect 408000 35000 433000 38000
rect 450000 37000 464000 39000
rect 482000 37000 495000 39000
rect 451000 35000 465000 37000
rect 481000 36000 495000 37000
rect 480000 35000 495000 36000
rect 409000 32000 432000 35000
rect 451000 34000 466000 35000
rect 480000 34000 494000 35000
rect 452000 33000 468000 34000
rect 478000 33000 494000 34000
rect 452000 32000 470000 33000
rect 477000 32000 493000 33000
rect 520000 32000 533000 79000
rect 566000 70000 579000 82000
rect 620000 70000 638000 71000
rect 675000 70000 689000 71000
rect 729000 70000 743000 71000
rect 554000 61000 597000 70000
rect 616000 69000 642000 70000
rect 672000 69000 706000 70000
rect 726000 69000 745000 70000
rect 613000 68000 644000 69000
rect 670000 68000 706000 69000
rect 724000 68000 747000 69000
rect 612000 67000 645000 68000
rect 668000 67000 706000 68000
rect 722000 67000 749000 68000
rect 612000 66000 646000 67000
rect 667000 66000 706000 67000
rect 721000 66000 750000 67000
rect 612000 65000 647000 66000
rect 666000 65000 706000 66000
rect 720000 65000 751000 66000
rect 612000 63000 648000 65000
rect 665000 63000 706000 65000
rect 719000 64000 752000 65000
rect 718000 63000 753000 64000
rect 612000 62000 649000 63000
rect 664000 62000 706000 63000
rect 612000 61000 624000 62000
rect 632000 61000 649000 62000
rect 566000 36000 579000 61000
rect 612000 60000 619000 61000
rect 634000 60000 649000 61000
rect 663000 61000 678000 62000
rect 685000 61000 706000 62000
rect 717000 62000 753000 63000
rect 717000 61000 733000 62000
rect 738000 61000 754000 62000
rect 663000 60000 676000 61000
rect 687000 60000 699000 61000
rect 716000 60000 730000 61000
rect 740000 60000 754000 61000
rect 612000 59000 616000 60000
rect 636000 59000 650000 60000
rect 612000 58000 614000 59000
rect 637000 56000 650000 59000
rect 663000 58000 675000 60000
rect 688000 58000 700000 60000
rect 716000 59000 729000 60000
rect 741000 59000 755000 60000
rect 715000 58000 728000 59000
rect 742000 58000 755000 59000
rect 638000 52000 650000 56000
rect 624000 51000 650000 52000
rect 620000 50000 650000 51000
rect 662000 51000 674000 58000
rect 689000 51000 701000 58000
rect 715000 57000 727000 58000
rect 714000 56000 727000 57000
rect 714000 53000 726000 56000
rect 743000 55000 756000 58000
rect 713000 52000 726000 53000
rect 744000 52000 756000 55000
rect 662000 50000 675000 51000
rect 617000 49000 650000 50000
rect 615000 48000 650000 49000
rect 614000 47000 650000 48000
rect 663000 49000 675000 50000
rect 688000 49000 700000 51000
rect 663000 48000 676000 49000
rect 687000 48000 700000 49000
rect 663000 47000 678000 48000
rect 685000 47000 700000 48000
rect 613000 46000 650000 47000
rect 664000 46000 699000 47000
rect 612000 45000 650000 46000
rect 611000 44000 650000 45000
rect 610000 43000 650000 44000
rect 610000 42000 627000 43000
rect 609000 41000 625000 42000
rect 609000 40000 623000 41000
rect 609000 39000 622000 40000
rect 608000 38000 622000 39000
rect 567000 34000 580000 36000
rect 608000 35000 621000 38000
rect 638000 37000 650000 43000
rect 665000 45000 699000 46000
rect 665000 44000 698000 45000
rect 665000 43000 697000 44000
rect 713000 43000 756000 52000
rect 665000 42000 696000 43000
rect 664000 41000 695000 42000
rect 663000 40000 693000 41000
rect 713000 40000 725000 43000
rect 663000 39000 691000 40000
rect 637000 36000 650000 37000
rect 662000 38000 674000 39000
rect 676000 38000 688000 39000
rect 713000 38000 726000 40000
rect 662000 37000 673000 38000
rect 713000 37000 727000 38000
rect 662000 36000 672000 37000
rect 714000 36000 727000 37000
rect 636000 35000 650000 36000
rect 608000 34000 622000 35000
rect 634000 34000 650000 35000
rect 567000 33000 581000 34000
rect 609000 33000 622000 34000
rect 633000 33000 650000 34000
rect 567000 32000 582000 33000
rect 596000 32000 597000 33000
rect 410000 31000 432000 32000
rect 453000 31000 493000 32000
rect 410000 29000 431000 31000
rect 453000 30000 492000 31000
rect 411000 28000 431000 29000
rect 454000 28000 491000 30000
rect 411000 26000 430000 28000
rect 455000 27000 490000 28000
rect 456000 26000 489000 27000
rect 412000 25000 430000 26000
rect 457000 25000 487000 26000
rect 412000 22000 429000 25000
rect 459000 24000 486000 25000
rect 461000 23000 484000 24000
rect 463000 22000 482000 23000
rect 505000 22000 547000 32000
rect 567000 31000 584000 32000
rect 591000 31000 597000 32000
rect 567000 30000 597000 31000
rect 568000 28000 597000 30000
rect 609000 32000 623000 33000
rect 632000 32000 650000 33000
rect 609000 31000 625000 32000
rect 630000 31000 650000 32000
rect 661000 34000 673000 36000
rect 714000 35000 728000 36000
rect 714000 34000 729000 35000
rect 661000 33000 674000 34000
rect 715000 33000 730000 34000
rect 661000 32000 676000 33000
rect 715000 32000 732000 33000
rect 750000 32000 754000 33000
rect 661000 31000 693000 32000
rect 716000 31000 735000 32000
rect 744000 31000 754000 32000
rect 609000 29000 650000 31000
rect 662000 30000 697000 31000
rect 716000 30000 754000 31000
rect 662000 29000 699000 30000
rect 717000 29000 754000 30000
rect 569000 26000 597000 28000
rect 610000 27000 650000 29000
rect 663000 28000 701000 29000
rect 663000 27000 702000 28000
rect 718000 27000 754000 29000
rect 611000 26000 638000 27000
rect 570000 25000 597000 26000
rect 612000 25000 637000 26000
rect 571000 24000 597000 25000
rect 613000 24000 636000 25000
rect 573000 23000 597000 24000
rect 614000 23000 634000 24000
rect 575000 22000 597000 23000
rect 616000 22000 632000 23000
rect 639000 22000 650000 27000
rect 664000 26000 703000 27000
rect 720000 26000 754000 27000
rect 665000 25000 704000 26000
rect 721000 25000 754000 26000
rect 664000 24000 704000 25000
rect 722000 24000 754000 25000
rect 662000 23000 705000 24000
rect 724000 23000 754000 24000
rect 662000 22000 676000 23000
rect 685000 22000 705000 23000
rect 726000 22000 750000 23000
rect 8000 21000 21000 22000
rect 54000 21000 64000 22000
rect 97000 21000 109000 22000
rect 242000 21000 256000 22000
rect 272000 21000 287000 22000
rect 467000 21000 478000 22000
rect 579000 21000 591000 22000
rect 619000 21000 628000 22000
rect 661000 21000 675000 22000
rect 690000 21000 705000 22000
rect 730000 21000 744000 22000
rect 8000 20000 20000 21000
rect 7000 19000 19000 20000
rect 6000 18000 19000 19000
rect 54000 19000 63000 21000
rect 97000 20000 110000 21000
rect 242000 20000 255000 21000
rect 273000 20000 287000 21000
rect 98000 19000 110000 20000
rect 54000 18000 62000 19000
rect 99000 18000 111000 19000
rect 241000 18000 254000 20000
rect 6000 17000 18000 18000
rect 54000 17000 61000 18000
rect 99000 17000 112000 18000
rect 5000 16000 18000 17000
rect 55000 16000 61000 17000
rect 100000 16000 112000 17000
rect 5000 15000 17000 16000
rect 4000 14000 17000 15000
rect 55000 15000 60000 16000
rect 100000 15000 113000 16000
rect 4000 13000 16000 14000
rect 55000 13000 59000 15000
rect 101000 14000 113000 15000
rect 241000 15000 253000 18000
rect 274000 16000 287000 20000
rect 660000 19000 673000 21000
rect 692000 19000 706000 21000
rect 273000 15000 287000 16000
rect 241000 14000 254000 15000
rect 273000 14000 286000 15000
rect 101000 13000 114000 14000
rect 3000 12000 15000 13000
rect 55000 12000 58000 13000
rect 102000 12000 114000 13000
rect 241000 13000 255000 14000
rect 272000 13000 286000 14000
rect 241000 12000 257000 13000
rect 269000 12000 286000 13000
rect 659000 14000 672000 19000
rect 693000 17000 706000 19000
rect 693000 16000 705000 17000
rect 692000 15000 705000 16000
rect 691000 14000 705000 15000
rect 659000 13000 673000 14000
rect 690000 13000 705000 14000
rect 659000 12000 675000 13000
rect 688000 12000 704000 13000
rect 2000 11000 15000 12000
rect 56000 11000 57000 12000
rect 103000 11000 115000 12000
rect 241000 11000 262000 12000
rect 264000 11000 285000 12000
rect 660000 11000 680000 12000
rect 683000 11000 704000 12000
rect 2000 10000 14000 11000
rect 103000 10000 116000 11000
rect 1000 9000 116000 10000
rect 242000 10000 284000 11000
rect 660000 10000 703000 11000
rect 242000 9000 283000 10000
rect 661000 9000 702000 10000
rect 1000 8000 117000 9000
rect 243000 8000 282000 9000
rect 661000 8000 701000 9000
rect 0 7000 117000 8000
rect 244000 7000 281000 8000
rect 662000 7000 700000 8000
rect 0 3000 118000 7000
rect 245000 6000 280000 7000
rect 664000 6000 698000 7000
rect 247000 5000 278000 6000
rect 665000 5000 697000 6000
rect 249000 4000 276000 5000
rect 668000 4000 694000 5000
rect 253000 3000 272000 4000
rect 671000 3000 691000 4000
rect 0 2000 117000 3000
rect 1000 1000 117000 2000
rect 1000 0 116000 1000
<< end >>
