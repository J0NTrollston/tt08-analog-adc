magic
tech sky130A
timestamp 1730258808
<< metal2 >>
rect 4560 4260 4670 4270
rect 5020 4260 5100 4270
rect 4540 4250 4700 4260
rect 5020 4250 5170 4260
rect 4520 4240 4720 4250
rect 5020 4240 5200 4250
rect 4500 4230 4730 4240
rect 5020 4230 5210 4240
rect 4490 4220 4740 4230
rect 5020 4220 5220 4230
rect 4480 4210 4606 4220
rect 4620 4210 4750 4220
rect 4470 4200 4570 4210
rect 4670 4200 4760 4210
rect 4470 4190 4550 4200
rect 4680 4190 4770 4200
rect 4460 4180 4540 4190
rect 4700 4180 4770 4190
rect 4460 4170 4530 4180
rect 4710 4170 4780 4180
rect 4450 4160 4520 4170
rect 4720 4160 4780 4170
rect 4450 4150 4510 4160
rect 4720 4150 4790 4160
rect 4440 4140 4510 4150
rect 4440 4050 4500 4140
rect 4730 4130 4790 4150
rect 4740 4060 4800 4130
rect 4440 4040 4510 4050
rect 4450 4030 4510 4040
rect 4730 4030 4790 4060
rect 4450 4010 4520 4030
rect 4720 4020 4790 4030
rect 4710 4010 4780 4020
rect 4460 4000 4530 4010
rect 4700 4000 4780 4010
rect 4460 3990 4550 4000
rect 4690 3990 4770 4000
rect 4470 3980 4560 3990
rect 4680 3980 4760 3990
rect 4480 3970 4590 3980
rect 4650 3970 4760 3980
rect 5020 3980 5070 4220
rect 5130 4210 5230 4220
rect 5160 4200 5240 4210
rect 5170 4190 5250 4200
rect 5180 4180 5250 4190
rect 5190 4170 5260 4180
rect 5200 4140 5260 4170
rect 5210 4120 5260 4140
rect 5210 4070 5270 4120
rect 5210 4060 5260 4070
rect 5200 4030 5260 4060
rect 5190 4020 5260 4030
rect 5190 4010 5250 4020
rect 5180 4000 5250 4010
rect 5170 3990 5240 4000
rect 5140 3980 5230 3990
rect 5020 3970 5230 3980
rect 4490 3960 4750 3970
rect 5020 3960 5210 3970
rect 4500 3950 4740 3960
rect 5020 3950 5200 3960
rect 4510 3940 4720 3950
rect 5020 3940 5180 3950
rect 4530 3930 4710 3940
rect 5020 3930 5140 3940
rect 4550 3920 4690 3930
rect 4570 2960 4670 3920
rect 3820 2950 4670 2960
rect 3800 2940 4670 2950
rect 3790 2920 4670 2940
rect 2580 2450 2620 2460
rect 2050 2440 2140 2450
rect 2540 2440 2660 2450
rect 2020 2430 2160 2440
rect 2510 2430 2690 2440
rect 2010 2420 2180 2430
rect 2500 2420 2700 2430
rect 1990 2410 2190 2420
rect 2480 2410 2720 2420
rect 1980 2400 2190 2410
rect 2470 2400 2730 2410
rect 1970 2390 2060 2400
rect 2130 2390 2180 2400
rect 2460 2390 2570 2400
rect 2620 2390 2740 2400
rect 1970 2380 2040 2390
rect 2150 2380 2174 2390
rect 2460 2380 2550 2390
rect 2650 2380 2740 2390
rect 1960 2370 2030 2380
rect 2160 2370 2174 2380
rect 2450 2370 2530 2380
rect 2670 2370 2750 2380
rect 1960 2360 2020 2370
rect 2440 2360 2520 2370
rect 2680 2360 2760 2370
rect 1950 2340 2010 2360
rect 2440 2350 2510 2360
rect 2690 2350 2760 2360
rect 2430 2340 2500 2350
rect 2700 2340 2770 2350
rect 1950 2330 2000 2340
rect 1940 2220 2000 2330
rect 2430 2320 2490 2340
rect 2710 2330 2770 2340
rect 3460 2330 3600 2920
rect 2710 2320 3440 2330
rect 3454 2320 3600 2330
rect 2080 2290 2104 2294
rect 2080 2280 2200 2290
rect 2090 2266 2200 2280
rect 2080 2250 2200 2266
rect 2090 2240 2104 2250
rect 1950 2200 2010 2220
rect 1950 2190 2020 2200
rect 1960 2180 2030 2190
rect 1960 2170 2040 2180
rect 2150 2170 2200 2250
rect 2420 2230 2480 2320
rect 2710 2310 3600 2320
rect 2720 2240 3600 2310
rect 2710 2230 3600 2240
rect 2430 2210 2490 2230
rect 2710 2210 2770 2230
rect 3450 2220 3600 2230
rect 2430 2200 2500 2210
rect 2700 2200 2770 2210
rect 2440 2190 2510 2200
rect 2690 2190 2760 2200
rect 2440 2180 2520 2190
rect 2680 2180 2760 2190
rect 2450 2170 2530 2180
rect 2670 2170 2750 2180
rect 1970 2160 2050 2170
rect 2140 2160 2200 2170
rect 1980 2150 2200 2160
rect 2460 2160 2550 2170
rect 2650 2160 2740 2170
rect 2460 2150 2580 2160
rect 2620 2150 2730 2160
rect 1990 2140 2200 2150
rect 2470 2140 2730 2150
rect 2000 2130 2190 2140
rect 2490 2130 2710 2140
rect 2020 2120 2170 2130
rect 2500 2120 2700 2130
rect 2040 2110 2150 2120
rect 2510 2110 2680 2120
rect 2540 2100 2660 2110
rect 2580 2090 2610 2100
rect 3460 1640 3600 2220
rect 3780 2890 4670 2920
rect 3780 2880 4660 2890
rect 3780 2870 4650 2880
rect 3780 2860 4640 2870
rect 3780 2284 3880 2860
rect 4240 2450 4260 2460
rect 5340 2450 5400 2460
rect 4230 2440 4260 2450
rect 5310 2440 5430 2450
rect 5770 2440 5890 2450
rect 4200 2430 4260 2440
rect 5280 2430 5450 2440
rect 5770 2430 5950 2440
rect 4180 2420 4260 2430
rect 5270 2420 5470 2430
rect 5770 2420 5960 2430
rect 4160 2410 4260 2420
rect 5250 2410 5490 2420
rect 4140 2400 4260 2410
rect 5240 2400 5500 2410
rect 5770 2400 5980 2420
rect 4130 2390 4260 2400
rect 4100 2380 4260 2390
rect 5230 2390 5340 2400
rect 5400 2390 5510 2400
rect 5230 2380 5320 2390
rect 5420 2380 5510 2390
rect 4080 2370 4260 2380
rect 5220 2370 5300 2380
rect 5440 2370 5520 2380
rect 4070 2360 4260 2370
rect 4040 2350 4260 2360
rect 5210 2360 5290 2370
rect 5450 2360 5530 2370
rect 5210 2350 5280 2360
rect 5460 2350 5530 2360
rect 4020 2340 4260 2350
rect 4000 2330 4260 2340
rect 5200 2340 5270 2350
rect 5470 2340 5540 2350
rect 5200 2330 5260 2340
rect 3990 2320 4260 2330
rect 4274 2320 5260 2330
rect 5480 2320 5540 2340
rect 3970 2310 5250 2320
rect 5480 2310 5550 2320
rect 3940 2300 5250 2310
rect 3920 2290 5250 2300
rect 3910 2284 5250 2290
rect 3780 2270 5250 2284
rect 3780 1690 3880 2270
rect 3910 2260 5250 2270
rect 3930 2250 5250 2260
rect 3950 2240 5250 2250
rect 5490 2240 5550 2310
rect 3970 2230 5250 2240
rect 5480 2230 5550 2240
rect 5770 2310 5830 2400
rect 5910 2390 5990 2400
rect 5930 2370 5990 2390
rect 5940 2340 5990 2370
rect 5930 2330 5990 2340
rect 5930 2320 5980 2330
rect 5910 2310 5980 2320
rect 5770 2300 5970 2310
rect 5770 2280 5950 2300
rect 5770 2270 5980 2280
rect 3990 2220 4260 2230
rect 4010 2210 4260 2220
rect 4030 2200 4260 2210
rect 5200 2210 5260 2230
rect 5480 2220 5540 2230
rect 5200 2200 5270 2210
rect 5470 2200 5540 2220
rect 4050 2190 4260 2200
rect 4070 2180 4260 2190
rect 5210 2190 5280 2200
rect 5460 2190 5530 2200
rect 5210 2180 5290 2190
rect 5450 2180 5530 2190
rect 4090 2170 4260 2180
rect 5220 2170 5300 2180
rect 5440 2170 5520 2180
rect 4110 2160 4260 2170
rect 4130 2150 4260 2160
rect 5230 2160 5320 2170
rect 5420 2160 5510 2170
rect 5770 2160 5830 2270
rect 5844 2260 5990 2270
rect 5930 2250 6000 2260
rect 5940 2240 6000 2250
rect 5950 2180 6010 2240
rect 5940 2170 6000 2180
rect 5920 2160 6000 2170
rect 5230 2150 5350 2160
rect 5390 2150 5500 2160
rect 4150 2140 4260 2150
rect 5240 2140 5500 2150
rect 5770 2140 5990 2160
rect 4170 2130 4260 2140
rect 5260 2130 5480 2140
rect 5770 2130 5970 2140
rect 4190 2120 4260 2130
rect 5270 2120 5470 2130
rect 5770 2120 5950 2130
rect 4210 2110 4260 2120
rect 5280 2110 5450 2120
rect 5770 2110 5920 2120
rect 4230 2100 4264 2110
rect 5310 2100 5430 2110
rect 4250 2090 4264 2100
rect 5360 2090 5380 2100
rect 3780 1680 4640 1690
rect 3780 1660 4660 1680
rect 3780 1640 4670 1660
rect 3790 1610 4670 1640
rect 3800 1600 4670 1610
rect 3820 1590 4670 1600
rect 4570 630 4670 1590
rect 5110 630 5160 640
rect 4550 620 4690 630
rect 5080 620 5200 630
rect 4530 610 4710 620
rect 5070 610 5220 620
rect 4510 600 4720 610
rect 5050 604 5230 610
rect 4500 590 4740 600
rect 5050 590 5240 604
rect 4490 580 4750 590
rect 5040 580 5120 590
rect 5160 580 5230 590
rect 4480 570 4580 580
rect 4650 570 4760 580
rect 4470 560 4560 570
rect 4680 560 4760 570
rect 5030 570 5100 580
rect 5190 570 5230 580
rect 4460 550 4540 560
rect 4690 550 4770 560
rect 4460 540 4530 550
rect 4700 540 4780 550
rect 4450 520 4520 540
rect 4710 530 4780 540
rect 5030 530 5090 570
rect 5200 560 5220 570
rect 4450 510 4510 520
rect 4720 510 4790 530
rect 5030 520 5100 530
rect 5030 510 5110 520
rect 4440 500 4510 510
rect 4730 500 4790 510
rect 5040 500 5130 510
rect 4440 410 4500 500
rect 4730 490 4800 500
rect 5040 490 5150 500
rect 4740 430 4800 490
rect 5050 480 5180 490
rect 5060 470 5200 480
rect 5080 460 5210 470
rect 5100 450 5230 460
rect 5120 440 5240 450
rect 5140 430 5240 440
rect 4730 420 4800 430
rect 5160 420 5250 430
rect 4440 400 4510 410
rect 4730 400 4790 420
rect 5180 410 5250 420
rect 4450 390 4510 400
rect 4720 390 4790 400
rect 4450 380 4520 390
rect 4720 380 4780 390
rect 4460 370 4530 380
rect 4710 370 4780 380
rect 5040 370 5054 380
rect 4460 360 4540 370
rect 4700 360 4770 370
rect 5040 360 5070 370
rect 5190 360 5250 410
rect 4470 350 4550 360
rect 4680 350 4770 360
rect 5030 350 5080 360
rect 5180 350 5250 360
rect 4480 340 4570 350
rect 4660 340 4760 350
rect 5020 340 5110 350
rect 5160 340 5240 350
rect 4480 330 4750 340
rect 5020 330 5230 340
rect 4500 320 4740 330
rect 5030 320 5230 330
rect 4510 310 4730 320
rect 5050 310 5210 320
rect 4520 300 4710 310
rect 5070 300 5200 310
rect 4540 290 4700 300
rect 5100 290 5170 300
rect 4560 280 4670 290
<< end >>
