** sch_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp_ladder_tb.sch
**.subckt opamp_ladder_tb out0 out1 out2 out3 in out0_parax out1_parax out2_parax out3_parax in
*.opin out0
*.opin out1
*.opin out2
*.opin out3
*.ipin in
*.opin out0_parax
*.opin out1_parax
*.opin out2_parax
*.opin out3_parax
*.ipin in
x1 VDD in VSS out3 out2 out1 out0 opamp_ladder
V1 VSS GND 0
V2 VDD GND 1.8
x2 in out3_parax out2_parax out1_parax out0_parax VSS VDD opamp_ladder_parax
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt





v_in in 0 1.8
.control
dc v_in 0 1.8 0.01
save all
write opamp_ladder_tb.raw
.endc



**** end user architecture code
**.ends

* expanding   symbol:  opamp_ladder.sym # of pins=7
** sym_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp_ladder.sym
** sch_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp_ladder.sch
.subckt opamp_ladder VDD in VSS out3 out2 out1 out0
*.opin out0
*.opin out2
*.opin out3
*.ipin in
*.iopin VDD
*.iopin VSS
*.opin out1
x1 VDD VSS node_0 in out0 VSS opamp
XR2 VSS node_0 VSS sky130_fd_pr__res_generic_nd W=1 L=8.4 mult=1 m=1
XR3 node_0 node_1 VSS sky130_fd_pr__res_generic_nd W=1 L=8.4 mult=1 m=1
XR4 node_1 node_2 VSS sky130_fd_pr__res_generic_nd W=1 L=8.4 mult=1 m=1
XR5 node_2 node_3 VSS sky130_fd_pr__res_generic_nd W=1 L=8.4 mult=1 m=1
x2 VDD VSS node_1 in out1 VSS opamp
x3 VDD VSS node_2 in out2 VSS opamp
x4 VDD VSS node_3 in out3 VSS opamp
XR1 node_3 VDD VSS sky130_fd_pr__res_generic_nd W=1 L=8.4 mult=1 m=1
.ends


* expanding   symbol:  opamp_ladder_parax.sym # of pins=7
** sym_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp_ladder.sym
.include /home/ttuser/Documents/tt08-analog-adc/mag/opamp_ladder.sim.spice

* expanding   symbol:  opamp.sym # of pins=6
** sym_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp.sym
** sch_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp.sch
.subckt opamp VDD ZREF vin_n vin_p Vout VGND
*.ipin vin_n
*.ipin vin_p
*.opin Vout
*.iopin VDD
*.iopin ZREF
*.iopin VGND
XM1 net1 vin_n net3 net3 sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 vin_p net3 net3 sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 net1 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 net1 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net3 VGND VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vout VGND VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 ZREF VGND VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net4 VDD net2 VGND sky130_fd_pr__nfet_01v8 L=0.6 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC1 net4 Vout sky130_fd_pr__cap_mim_m3_1 W=17.55 L=15 MF=1 m=1
XM6 Vout net2 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR1 ZREF VDD VGND sky130_fd_pr__res_generic_nd W=1 L=5 mult=1 m=1
XR2 VGND ZREF VGND sky130_fd_pr__res_generic_nd W=1 L=5 mult=1 m=1
.ends

.GLOBAL GND
.end
