magic
tech sky130A
timestamp 1730256539
<< metal2 >>
rect 5180 11130 6020 11200
rect 4620 11060 6580 11130
rect 4270 10990 6930 11060
rect 3990 10920 7210 10990
rect 3780 10850 7420 10920
rect 3570 10780 7630 10850
rect 3430 10710 7770 10780
rect 3290 10640 7910 10710
rect 3150 10570 8050 10640
rect 3010 10500 8260 10570
rect 2870 10430 8330 10500
rect 2730 10360 8470 10430
rect 2590 10290 8610 10360
rect 2520 10220 8680 10290
rect 2380 10150 8820 10220
rect 2310 10080 8890 10150
rect 2240 10010 8960 10080
rect 2100 9940 9100 10010
rect 2030 9870 9170 9940
rect 1960 9800 9240 9870
rect 1890 9730 9310 9800
rect 6370 9660 8470 9730
rect 8540 9660 9380 9730
rect 6370 9590 8400 9660
rect 6300 9450 8400 9590
rect 8540 9590 9450 9660
rect 8540 9520 9520 9590
rect 8540 9450 9590 9520
rect 6230 9310 8330 9450
rect 8610 9380 9660 9450
rect 8610 9310 9730 9380
rect 6160 9240 8260 9310
rect 8610 9240 9800 9310
rect 6160 9170 8190 9240
rect 6090 9100 8190 9170
rect 8610 9170 9870 9240
rect 8610 9100 9940 9170
rect 6090 9030 8120 9100
rect 6020 8960 8120 9030
rect 8680 8960 10010 9100
rect 6020 8890 8050 8960
rect 5950 8820 8050 8890
rect 8680 8890 10080 8960
rect 8680 8820 10150 8890
rect 5950 8750 7980 8820
rect 5880 8680 7980 8750
rect 8750 8680 10220 8820
rect 5880 8610 7910 8680
rect 5810 8540 7910 8610
rect 8750 8610 10290 8680
rect 5810 8470 7840 8540
rect 8750 8470 10360 8610
rect 5740 8400 7840 8470
rect 770 8330 4270 8400
rect 5740 8330 7770 8400
rect 700 8260 4270 8330
rect 5670 8260 7770 8330
rect 8820 8330 10430 8470
rect 630 8120 4200 8260
rect 5600 8120 7700 8260
rect 8820 8190 10500 8330
rect 560 7980 4130 8120
rect 5600 8050 7630 8120
rect 5530 7980 7630 8050
rect 8890 8050 10570 8190
rect 560 7910 4060 7980
rect 5530 7910 7560 7980
rect 490 7840 4060 7910
rect 5460 7840 7560 7910
rect 8890 7910 10640 8050
rect 8890 7840 10710 7910
rect 490 7770 3990 7840
rect 420 7700 3990 7770
rect 5390 7700 7490 7840
rect 8960 7770 10710 7840
rect 420 7630 3920 7700
rect 350 7560 3920 7630
rect 5320 7560 7420 7700
rect 8960 7630 10780 7770
rect 350 7420 3850 7560
rect 5250 7420 7350 7560
rect 8960 7490 10850 7630
rect 9030 7420 10850 7490
rect 280 7280 3780 7420
rect 5180 7280 7280 7420
rect 280 7210 3710 7280
rect 210 7140 3710 7210
rect 5110 7140 7210 7280
rect 9030 7210 10920 7420
rect 210 7000 3640 7140
rect 5040 7000 7140 7140
rect 210 6930 3570 7000
rect 140 6860 3570 6930
rect 4970 6860 7070 7000
rect 9100 6930 10990 7210
rect 9100 6860 11060 6930
rect 140 6720 3500 6860
rect 4900 6720 7000 6860
rect 140 6580 3430 6720
rect 4830 6580 6930 6720
rect 9170 6580 11060 6860
rect 70 6440 3360 6580
rect 4760 6440 6860 6580
rect 9170 6510 11130 6580
rect 70 6300 3290 6440
rect 4690 6300 6790 6440
rect 70 6160 3220 6300
rect 4620 6160 6720 6300
rect 9240 6230 11130 6510
rect 70 6020 3150 6160
rect 4550 6020 6650 6160
rect 7980 6090 8050 6160
rect 7980 6020 8120 6090
rect 0 5880 3080 6020
rect 4480 5880 6580 6020
rect 7910 5880 8120 6020
rect 9310 6020 11130 6230
rect 9310 5880 11200 6020
rect 0 5740 3010 5880
rect 4410 5740 6510 5880
rect 7840 5740 8120 5880
rect 0 5600 2940 5740
rect 4340 5600 6440 5740
rect 7770 5600 8190 5740
rect 0 5460 2870 5600
rect 4270 5460 6370 5600
rect 7700 5460 8190 5600
rect 9380 5530 11200 5880
rect 0 5320 2800 5460
rect 4200 5320 6300 5460
rect 7630 5320 8260 5460
rect 0 5180 2730 5320
rect 4130 5180 6230 5320
rect 7560 5180 8260 5320
rect 9450 5250 11200 5530
rect 70 5040 2660 5180
rect 4060 5040 6160 5180
rect 7490 5110 8260 5180
rect 9520 5180 11200 5250
rect 7490 5040 8330 5110
rect 70 4900 2590 5040
rect 3990 4900 6090 5040
rect 7420 4900 8330 5040
rect 9520 4900 11130 5180
rect 70 4760 2520 4900
rect 3920 4760 6020 4900
rect 7350 4830 8330 4900
rect 7350 4760 8400 4830
rect 70 4620 2450 4760
rect 3850 4620 5950 4760
rect 7280 4620 8400 4760
rect 140 4480 2380 4620
rect 3780 4480 5880 4620
rect 7210 4480 8400 4620
rect 9590 4620 11130 4900
rect 9590 4550 11060 4620
rect 140 4340 2310 4480
rect 3710 4410 4760 4480
rect 4900 4410 5810 4480
rect 3710 4340 4690 4410
rect 5110 4340 5810 4410
rect 7140 4340 8470 4480
rect 140 4270 2240 4340
rect 210 4200 2240 4270
rect 3640 4270 4690 4340
rect 5320 4270 5740 4340
rect 3640 4200 4620 4270
rect 5530 4200 5740 4270
rect 7070 4200 8470 4340
rect 9660 4270 11060 4550
rect 210 4060 2170 4200
rect 3570 4130 4620 4200
rect 7000 4130 8470 4200
rect 3570 4060 4550 4130
rect 7000 4060 8540 4130
rect 210 3990 2100 4060
rect 3500 3990 4550 4060
rect 280 3920 2100 3990
rect 6930 3920 8540 4060
rect 9730 3990 10990 4270
rect 9730 3920 10920 3990
rect 280 3780 2030 3920
rect 6860 3850 8540 3920
rect 6860 3780 8610 3850
rect 350 3640 1960 3780
rect 6930 3710 8610 3780
rect 7140 3640 8610 3710
rect 350 3570 1890 3640
rect 7350 3570 8610 3640
rect 9800 3780 10920 3920
rect 9800 3570 10850 3780
rect 420 3500 1890 3570
rect 7560 3500 8610 3570
rect 420 3430 1820 3500
rect 7770 3430 8680 3500
rect 490 3360 1820 3430
rect 7980 3360 8680 3430
rect 490 3290 1750 3360
rect 560 3220 1750 3290
rect 8190 3220 8680 3360
rect 9870 3430 10780 3570
rect 9870 3290 10710 3430
rect 560 3150 1680 3220
rect 7980 3150 8680 3220
rect 9940 3150 10640 3290
rect 630 3010 1610 3150
rect 7700 3080 8750 3150
rect 7420 3010 8750 3080
rect 700 2940 1610 3010
rect 7140 2940 8750 3010
rect 9940 3010 10570 3150
rect 9940 2940 10500 3010
rect 700 2870 1540 2940
rect 6860 2870 8750 2940
rect 10010 2870 10500 2940
rect 770 2800 1540 2870
rect 6650 2800 8820 2870
rect 770 2730 1470 2800
rect 6370 2730 8820 2800
rect 840 2660 1470 2730
rect 6090 2660 8820 2730
rect 10010 2730 10430 2870
rect 10010 2660 10360 2730
rect 840 2590 3850 2660
rect 5810 2590 8820 2660
rect 910 2520 3780 2590
rect 5530 2520 8820 2590
rect 10080 2590 10360 2660
rect 10080 2520 10290 2590
rect 980 2450 3780 2520
rect 5250 2450 6020 2520
rect 980 2380 3710 2450
rect 4970 2380 5810 2450
rect 6160 2380 8890 2520
rect 1050 2310 3710 2380
rect 4760 2310 5670 2380
rect 1120 2240 3640 2310
rect 4480 2240 5460 2310
rect 6090 2240 8890 2380
rect 10080 2380 10220 2520
rect 10080 2310 10150 2380
rect 1190 2170 3640 2240
rect 4200 2170 5320 2240
rect 1190 2100 3570 2170
rect 3920 2100 5110 2170
rect 6020 2100 8960 2240
rect 1260 2030 3570 2100
rect 3640 2030 4970 2100
rect 1330 1960 4760 2030
rect 5950 1960 8960 2100
rect 1400 1890 4620 1960
rect 5880 1890 8960 1960
rect 1470 1820 4550 1890
rect 5880 1820 9030 1890
rect 1540 1750 4480 1820
rect 1610 1680 4480 1750
rect 5810 1680 9030 1820
rect 1680 1610 4410 1680
rect 1750 1540 4410 1610
rect 5740 1540 9030 1680
rect 1820 1470 4340 1540
rect 1890 1400 4340 1470
rect 5670 1400 9100 1540
rect 1960 1330 4270 1400
rect 2030 1260 4270 1330
rect 5600 1260 9100 1400
rect 2100 1190 4200 1260
rect 2240 1120 4200 1190
rect 5530 1190 9100 1260
rect 5530 1120 8960 1190
rect 2310 1050 4130 1120
rect 2380 980 4130 1050
rect 5460 1050 8890 1120
rect 5460 980 8820 1050
rect 2520 910 4060 980
rect 2590 840 4060 910
rect 5390 910 8680 980
rect 5390 840 8610 910
rect 2730 770 3990 840
rect 2870 700 3990 770
rect 5320 770 8470 840
rect 5320 700 8330 770
rect 3010 630 3920 700
rect 3150 560 3920 630
rect 5250 630 8190 700
rect 5250 560 8050 630
rect 3290 490 3850 560
rect 5180 490 7910 560
rect 3430 420 3850 490
rect 5110 420 7770 490
rect 3570 350 3780 420
rect 5110 350 7630 420
rect 5040 280 7420 350
rect 5040 210 7210 280
rect 5040 140 6930 210
rect 4970 70 6580 140
rect 5180 0 6020 70
<< end >>
