magic
tech sky130A
magscale 1 2
timestamp 1730221101
<< viali >>
rect 9321 9129 9355 9163
rect 9137 8993 9171 9027
rect 8585 8925 8619 8959
rect 9045 8925 9079 8959
rect 8953 8857 8987 8891
rect 10425 8585 10459 8619
rect 10701 8585 10735 8619
rect 3341 8381 3375 8415
rect 5365 8381 5399 8415
rect 7481 8381 7515 8415
rect 7941 8381 7975 8415
rect 8125 8381 8159 8415
rect 8585 8381 8619 8415
rect 8861 8381 8895 8415
rect 9045 8381 9079 8415
rect 10517 8381 10551 8415
rect 3608 8313 3642 8347
rect 5632 8313 5666 8347
rect 6837 8313 6871 8347
rect 9290 8313 9324 8347
rect 4721 8245 4755 8279
rect 6745 8245 6779 8279
rect 8401 8245 8435 8279
rect 8769 8245 8803 8279
rect 3525 8041 3559 8075
rect 4261 8041 4295 8075
rect 8493 8041 8527 8075
rect 3709 7973 3743 8007
rect 5181 7973 5215 8007
rect 3249 7905 3283 7939
rect 4169 7905 4203 7939
rect 4445 7905 4479 7939
rect 5365 7905 5399 7939
rect 6101 7905 6135 7939
rect 7205 7905 7239 7939
rect 9229 7905 9263 7939
rect 9485 7905 9519 7939
rect 5641 7837 5675 7871
rect 5917 7837 5951 7871
rect 6377 7837 6411 7871
rect 6469 7837 6503 7871
rect 3433 7769 3467 7803
rect 4077 7769 4111 7803
rect 5549 7769 5583 7803
rect 3709 7701 3743 7735
rect 4629 7701 4663 7735
rect 6285 7701 6319 7735
rect 7113 7701 7147 7735
rect 10609 7701 10643 7735
rect 3985 7497 4019 7531
rect 4169 7497 4203 7531
rect 6193 7497 6227 7531
rect 6561 7497 6595 7531
rect 7573 7497 7607 7531
rect 9045 7497 9079 7531
rect 3065 7429 3099 7463
rect 3801 7361 3835 7395
rect 4813 7361 4847 7395
rect 6929 7361 6963 7395
rect 7021 7361 7055 7395
rect 10609 7361 10643 7395
rect 1685 7293 1719 7327
rect 4629 7293 4663 7327
rect 6745 7293 6779 7327
rect 6837 7293 6871 7327
rect 7481 7293 7515 7327
rect 7849 7293 7883 7327
rect 7941 7293 7975 7327
rect 8033 7293 8067 7327
rect 8217 7293 8251 7327
rect 8401 7293 8435 7327
rect 8585 7293 8619 7327
rect 8677 7293 8711 7327
rect 8769 7293 8803 7327
rect 9321 7293 9355 7327
rect 9597 7293 9631 7327
rect 11069 7293 11103 7327
rect 1952 7225 1986 7259
rect 4137 7225 4171 7259
rect 4353 7225 4387 7259
rect 5058 7225 5092 7259
rect 7389 7225 7423 7259
rect 9137 7225 9171 7259
rect 10057 7225 10091 7259
rect 3249 7157 3283 7191
rect 4537 7157 4571 7191
rect 9505 7157 9539 7191
rect 10885 7157 10919 7191
rect 2329 6953 2363 6987
rect 3433 6953 3467 6987
rect 8125 6953 8159 6987
rect 1593 6817 1627 6851
rect 2513 6817 2547 6851
rect 2789 6817 2823 6851
rect 3249 6817 3283 6851
rect 3525 6817 3559 6851
rect 4169 6817 4203 6851
rect 4353 6817 4387 6851
rect 4537 6817 4571 6851
rect 7665 6817 7699 6851
rect 8217 6817 8251 6851
rect 9689 6817 9723 6851
rect 9873 6817 9907 6851
rect 10425 6817 10459 6851
rect 1777 6749 1811 6783
rect 1869 6749 1903 6783
rect 1961 6749 1995 6783
rect 2053 6749 2087 6783
rect 2697 6749 2731 6783
rect 5825 6749 5859 6783
rect 6193 6749 6227 6783
rect 3249 6681 3283 6715
rect 10241 6681 10275 6715
rect 1409 6613 1443 6647
rect 2237 6613 2271 6647
rect 3985 6613 4019 6647
rect 4445 6613 4479 6647
rect 7849 6613 7883 6647
rect 8309 6613 8343 6647
rect 9781 6613 9815 6647
rect 2697 6409 2731 6443
rect 5273 6409 5307 6443
rect 6285 6409 6319 6443
rect 7665 6409 7699 6443
rect 2421 6341 2455 6375
rect 2513 6341 2547 6375
rect 3065 6341 3099 6375
rect 1041 6205 1075 6239
rect 1308 6205 1342 6239
rect 5089 6205 5123 6239
rect 5181 6205 5215 6239
rect 5365 6205 5399 6239
rect 5457 6205 5491 6239
rect 5641 6205 5675 6239
rect 7849 6205 7883 6239
rect 8125 6205 8159 6239
rect 8585 6205 8619 6239
rect 8953 6205 8987 6239
rect 10425 6205 10459 6239
rect 3525 6137 3559 6171
rect 7573 6137 7607 6171
rect 2697 6069 2731 6103
rect 5641 6069 5675 6103
rect 8033 6069 8067 6103
rect 10985 6069 11019 6103
rect 2513 5865 2547 5899
rect 2697 5865 2731 5899
rect 2881 5865 2915 5899
rect 4905 5865 4939 5899
rect 6561 5865 6595 5899
rect 7113 5865 7147 5899
rect 7573 5865 7607 5899
rect 8033 5865 8067 5899
rect 8309 5865 8343 5899
rect 2329 5797 2363 5831
rect 3792 5797 3826 5831
rect 5365 5797 5399 5831
rect 2605 5729 2639 5763
rect 2973 5729 3007 5763
rect 5181 5729 5215 5763
rect 5457 5729 5491 5763
rect 5641 5729 5675 5763
rect 6745 5729 6779 5763
rect 7481 5729 7515 5763
rect 7941 5729 7975 5763
rect 8125 5729 8159 5763
rect 8217 5729 8251 5763
rect 9505 5729 9539 5763
rect 9689 5729 9723 5763
rect 1409 5661 1443 5695
rect 3249 5661 3283 5695
rect 3525 5661 3559 5695
rect 7757 5661 7791 5695
rect 3065 5593 3099 5627
rect 2053 5525 2087 5559
rect 3157 5525 3191 5559
rect 4997 5525 5031 5559
rect 5549 5525 5583 5559
rect 9597 5525 9631 5559
rect 4077 5321 4111 5355
rect 4261 5321 4295 5355
rect 8125 5321 8159 5355
rect 10793 5321 10827 5355
rect 1501 5253 1535 5287
rect 3249 5253 3283 5287
rect 2145 5185 2179 5219
rect 2329 5185 2363 5219
rect 4721 5185 4755 5219
rect 5089 5185 5123 5219
rect 8493 5185 8527 5219
rect 1225 5117 1259 5151
rect 1317 5117 1351 5151
rect 3249 5117 3283 5151
rect 3525 5117 3559 5151
rect 6561 5117 6595 5151
rect 7113 5117 7147 5151
rect 7297 5117 7331 5151
rect 7573 5117 7607 5151
rect 7752 5117 7786 5151
rect 7941 5117 7975 5151
rect 8861 5117 8895 5151
rect 10333 5117 10367 5151
rect 1501 5049 1535 5083
rect 2973 5049 3007 5083
rect 4445 5049 4479 5083
rect 7849 5049 7883 5083
rect 8125 5049 8159 5083
rect 1593 4981 1627 5015
rect 3433 4981 3467 5015
rect 4245 4981 4279 5015
rect 6745 4981 6779 5015
rect 7021 4981 7055 5015
rect 7481 4981 7515 5015
rect 10517 4981 10551 5015
rect 1133 4777 1167 4811
rect 2697 4777 2731 4811
rect 2789 4777 2823 4811
rect 6285 4777 6319 4811
rect 6929 4777 6963 4811
rect 8493 4777 8527 4811
rect 1584 4709 1618 4743
rect 8861 4709 8895 4743
rect 1041 4641 1075 4675
rect 1225 4641 1259 4675
rect 3709 4641 3743 4675
rect 3893 4641 3927 4675
rect 6285 4641 6319 4675
rect 6469 4641 6503 4675
rect 6837 4641 6871 4675
rect 8953 4641 8987 4675
rect 1317 4573 1351 4607
rect 3341 4573 3375 4607
rect 3525 4573 3559 4607
rect 3801 4573 3835 4607
rect 3985 4573 4019 4607
rect 9045 4573 9079 4607
rect 1685 4233 1719 4267
rect 7113 4233 7147 4267
rect 9781 4233 9815 4267
rect 7665 4165 7699 4199
rect 8401 4097 8435 4131
rect 9505 4097 9539 4131
rect 9597 4097 9631 4131
rect 2798 4029 2832 4063
rect 3065 4029 3099 4063
rect 4721 4029 4755 4063
rect 5917 4029 5951 4063
rect 6101 4029 6135 4063
rect 7297 4029 7331 4063
rect 7573 4029 7607 4063
rect 7849 4029 7883 4063
rect 8125 4029 8159 4063
rect 8585 4029 8619 4063
rect 8677 4029 8711 4063
rect 8861 4029 8895 4063
rect 9045 4029 9079 4063
rect 9137 4029 9171 4063
rect 9229 4029 9263 4063
rect 9873 4029 9907 4063
rect 7481 3961 7515 3995
rect 8401 3961 8435 3995
rect 9597 3961 9631 3995
rect 4813 3893 4847 3927
rect 6009 3893 6043 3927
rect 8033 3893 8067 3927
rect 3709 3689 3743 3723
rect 8493 3689 8527 3723
rect 9137 3689 9171 3723
rect 6377 3621 6411 3655
rect 8401 3621 8435 3655
rect 2329 3553 2363 3587
rect 2596 3553 2630 3587
rect 6009 3553 6043 3587
rect 6285 3553 6319 3587
rect 6653 3553 6687 3587
rect 7757 3553 7791 3587
rect 7941 3553 7975 3587
rect 8125 3553 8159 3587
rect 8677 3553 8711 3587
rect 8953 3553 8987 3587
rect 9321 3553 9355 3587
rect 9505 3553 9539 3587
rect 9597 3553 9631 3587
rect 10241 3553 10275 3587
rect 6377 3485 6411 3519
rect 7849 3485 7883 3519
rect 8401 3485 8435 3519
rect 8769 3485 8803 3519
rect 8861 3485 8895 3519
rect 10333 3485 10367 3519
rect 6193 3417 6227 3451
rect 6561 3417 6595 3451
rect 8217 3417 8251 3451
rect 9873 3417 9907 3451
rect 5825 3349 5859 3383
rect 2697 3145 2731 3179
rect 3249 3145 3283 3179
rect 8401 3145 8435 3179
rect 9045 3145 9079 3179
rect 9689 3145 9723 3179
rect 9873 3145 9907 3179
rect 10425 3145 10459 3179
rect 9597 3077 9631 3111
rect 3801 3009 3835 3043
rect 4905 3009 4939 3043
rect 6377 3009 6411 3043
rect 8125 3009 8159 3043
rect 8677 3009 8711 3043
rect 2697 2941 2731 2975
rect 2881 2941 2915 2975
rect 4629 2941 4663 2975
rect 8033 2941 8067 2975
rect 8585 2941 8619 2975
rect 8769 2941 8803 2975
rect 8861 2941 8895 2975
rect 9229 2941 9263 2975
rect 9873 2941 9907 2975
rect 10241 2941 10275 2975
rect 10333 2941 10367 2975
rect 10517 2941 10551 2975
rect 9321 2873 9355 2907
rect 9413 2805 9447 2839
rect 9045 2601 9079 2635
rect 9289 2533 9323 2567
rect 9505 2533 9539 2567
rect 5089 2465 5123 2499
rect 6009 2465 6043 2499
rect 6193 2465 6227 2499
rect 5181 2397 5215 2431
rect 8585 2397 8619 2431
rect 8953 2329 8987 2363
rect 5365 2261 5399 2295
rect 6193 2261 6227 2295
rect 9137 2261 9171 2295
rect 9321 2261 9355 2295
rect 2421 2057 2455 2091
rect 3801 2057 3835 2091
rect 6837 2057 6871 2091
rect 8769 2057 8803 2091
rect 5089 1921 5123 1955
rect 5365 1921 5399 1955
rect 7021 1853 7055 1887
rect 7205 1853 7239 1887
rect 8861 1853 8895 1887
rect 2697 1785 2731 1819
rect 3709 1785 3743 1819
rect 7113 1717 7147 1751
rect 8401 1717 8435 1751
rect 2697 1513 2731 1547
rect 2865 1513 2899 1547
rect 3525 1513 3559 1547
rect 3617 1513 3651 1547
rect 7665 1513 7699 1547
rect 10149 1513 10183 1547
rect 3065 1445 3099 1479
rect 3157 1445 3191 1479
rect 3357 1445 3391 1479
rect 3985 1377 4019 1411
rect 8217 1377 8251 1411
rect 10333 1377 10367 1411
rect 4077 1309 4111 1343
rect 5917 1309 5951 1343
rect 6193 1309 6227 1343
rect 8125 1309 8159 1343
rect 7849 1241 7883 1275
rect 2881 1173 2915 1207
rect 3341 1173 3375 1207
rect 1409 969 1443 1003
rect 3617 969 3651 1003
rect 6009 969 6043 1003
rect 8401 901 8435 935
rect 1225 765 1259 799
rect 3801 765 3835 799
rect 6193 765 6227 799
rect 8585 765 8619 799
<< metal1 >>
rect 552 9274 11568 9296
rect 552 9222 3112 9274
rect 3164 9222 3176 9274
rect 3228 9222 3240 9274
rect 3292 9222 3304 9274
rect 3356 9222 3368 9274
rect 3420 9222 5826 9274
rect 5878 9222 5890 9274
rect 5942 9222 5954 9274
rect 6006 9222 6018 9274
rect 6070 9222 6082 9274
rect 6134 9222 8540 9274
rect 8592 9222 8604 9274
rect 8656 9222 8668 9274
rect 8720 9222 8732 9274
rect 8784 9222 8796 9274
rect 8848 9222 11254 9274
rect 11306 9222 11318 9274
rect 11370 9222 11382 9274
rect 11434 9222 11446 9274
rect 11498 9222 11510 9274
rect 11562 9222 11568 9274
rect 552 9200 11568 9222
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 9309 9163 9367 9169
rect 9309 9160 9321 9163
rect 8352 9132 9321 9160
rect 8352 9120 8358 9132
rect 9309 9129 9321 9132
rect 9355 9129 9367 9163
rect 9309 9123 9367 9129
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 8993 9183 9027
rect 9125 8987 9183 8993
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 8662 8956 8668 8968
rect 8619 8928 8668 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 8662 8916 8668 8928
rect 8720 8916 8726 8968
rect 9033 8959 9091 8965
rect 9033 8925 9045 8959
rect 9079 8956 9091 8959
rect 9140 8956 9168 8987
rect 9079 8928 9168 8956
rect 9079 8925 9091 8928
rect 9033 8919 9091 8925
rect 8938 8848 8944 8900
rect 8996 8848 9002 8900
rect 552 8730 11408 8752
rect 552 8678 1755 8730
rect 1807 8678 1819 8730
rect 1871 8678 1883 8730
rect 1935 8678 1947 8730
rect 1999 8678 2011 8730
rect 2063 8678 4469 8730
rect 4521 8678 4533 8730
rect 4585 8678 4597 8730
rect 4649 8678 4661 8730
rect 4713 8678 4725 8730
rect 4777 8678 7183 8730
rect 7235 8678 7247 8730
rect 7299 8678 7311 8730
rect 7363 8678 7375 8730
rect 7427 8678 7439 8730
rect 7491 8678 9897 8730
rect 9949 8678 9961 8730
rect 10013 8678 10025 8730
rect 10077 8678 10089 8730
rect 10141 8678 10153 8730
rect 10205 8678 11408 8730
rect 552 8656 11408 8678
rect 8570 8576 8576 8628
rect 8628 8616 8634 8628
rect 8938 8616 8944 8628
rect 8628 8588 8944 8616
rect 8628 8576 8634 8588
rect 8938 8576 8944 8588
rect 8996 8616 9002 8628
rect 9398 8616 9404 8628
rect 8996 8588 9404 8616
rect 8996 8576 9002 8588
rect 9398 8576 9404 8588
rect 9456 8616 9462 8628
rect 10413 8619 10471 8625
rect 10413 8616 10425 8619
rect 9456 8588 10425 8616
rect 9456 8576 9462 8588
rect 10413 8585 10425 8588
rect 10459 8585 10471 8619
rect 10413 8579 10471 8585
rect 10686 8576 10692 8628
rect 10744 8576 10750 8628
rect 6730 8508 6736 8560
rect 6788 8548 6794 8560
rect 6788 8520 6914 8548
rect 6788 8508 6794 8520
rect 6886 8480 6914 8520
rect 8662 8480 8668 8492
rect 6886 8452 8668 8480
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8412 3387 8415
rect 3418 8412 3424 8424
rect 3375 8384 3424 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 4798 8372 4804 8424
rect 4856 8412 4862 8424
rect 7484 8421 7512 8452
rect 8662 8440 8668 8452
rect 8720 8480 8726 8492
rect 8720 8452 9168 8480
rect 8720 8440 8726 8452
rect 5353 8415 5411 8421
rect 5353 8412 5365 8415
rect 4856 8384 5365 8412
rect 4856 8372 4862 8384
rect 5353 8381 5365 8384
rect 5399 8381 5411 8415
rect 5353 8375 5411 8381
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8381 7527 8415
rect 7469 8375 7527 8381
rect 7929 8415 7987 8421
rect 7929 8381 7941 8415
rect 7975 8381 7987 8415
rect 7929 8375 7987 8381
rect 3602 8353 3608 8356
rect 3596 8307 3608 8353
rect 3602 8304 3608 8307
rect 3660 8304 3666 8356
rect 5626 8353 5632 8356
rect 5620 8307 5632 8353
rect 5626 8304 5632 8307
rect 5684 8304 5690 8356
rect 6825 8347 6883 8353
rect 6825 8344 6837 8347
rect 6656 8316 6837 8344
rect 4706 8236 4712 8288
rect 4764 8236 4770 8288
rect 6178 8236 6184 8288
rect 6236 8276 6242 8288
rect 6656 8276 6684 8316
rect 6825 8313 6837 8316
rect 6871 8313 6883 8347
rect 7944 8344 7972 8375
rect 8110 8372 8116 8424
rect 8168 8372 8174 8424
rect 8570 8372 8576 8424
rect 8628 8372 8634 8424
rect 8864 8421 8892 8452
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8381 8907 8415
rect 8849 8375 8907 8381
rect 9030 8372 9036 8424
rect 9088 8372 9094 8424
rect 9140 8412 9168 8452
rect 10505 8415 10563 8421
rect 10505 8412 10517 8415
rect 9140 8384 10517 8412
rect 10505 8381 10517 8384
rect 10551 8381 10563 8415
rect 10505 8375 10563 8381
rect 8588 8344 8616 8372
rect 7944 8316 8616 8344
rect 6825 8307 6883 8313
rect 8938 8304 8944 8356
rect 8996 8344 9002 8356
rect 9278 8347 9336 8353
rect 9278 8344 9290 8347
rect 8996 8316 9290 8344
rect 8996 8304 9002 8316
rect 9278 8313 9290 8316
rect 9324 8313 9336 8347
rect 9278 8307 9336 8313
rect 6236 8248 6684 8276
rect 6236 8236 6242 8248
rect 6730 8236 6736 8288
rect 6788 8236 6794 8288
rect 8294 8236 8300 8288
rect 8352 8276 8358 8288
rect 8389 8279 8447 8285
rect 8389 8276 8401 8279
rect 8352 8248 8401 8276
rect 8352 8236 8358 8248
rect 8389 8245 8401 8248
rect 8435 8245 8447 8279
rect 8389 8239 8447 8245
rect 8757 8279 8815 8285
rect 8757 8245 8769 8279
rect 8803 8276 8815 8279
rect 9122 8276 9128 8288
rect 8803 8248 9128 8276
rect 8803 8245 8815 8248
rect 8757 8239 8815 8245
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 552 8186 11568 8208
rect 552 8134 3112 8186
rect 3164 8134 3176 8186
rect 3228 8134 3240 8186
rect 3292 8134 3304 8186
rect 3356 8134 3368 8186
rect 3420 8134 5826 8186
rect 5878 8134 5890 8186
rect 5942 8134 5954 8186
rect 6006 8134 6018 8186
rect 6070 8134 6082 8186
rect 6134 8134 8540 8186
rect 8592 8134 8604 8186
rect 8656 8134 8668 8186
rect 8720 8134 8732 8186
rect 8784 8134 8796 8186
rect 8848 8134 11254 8186
rect 11306 8134 11318 8186
rect 11370 8134 11382 8186
rect 11434 8134 11446 8186
rect 11498 8134 11510 8186
rect 11562 8134 11568 8186
rect 552 8112 11568 8134
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8041 3571 8075
rect 3513 8035 3571 8041
rect 3237 7939 3295 7945
rect 3237 7905 3249 7939
rect 3283 7936 3295 7939
rect 3528 7936 3556 8035
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 4212 8044 4261 8072
rect 4212 8032 4218 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 4249 8035 4307 8041
rect 4798 8032 4804 8084
rect 4856 8072 4862 8084
rect 8481 8075 8539 8081
rect 8481 8072 8493 8075
rect 4856 8044 8493 8072
rect 4856 8032 4862 8044
rect 8481 8041 8493 8044
rect 8527 8041 8539 8075
rect 8481 8035 8539 8041
rect 3697 8007 3755 8013
rect 3697 7973 3709 8007
rect 3743 8004 3755 8007
rect 5169 8007 5227 8013
rect 3743 7976 5120 8004
rect 3743 7973 3755 7976
rect 3697 7967 3755 7973
rect 3283 7908 3556 7936
rect 3283 7905 3295 7908
rect 3237 7899 3295 7905
rect 3970 7896 3976 7948
rect 4028 7936 4034 7948
rect 4157 7939 4215 7945
rect 4157 7936 4169 7939
rect 4028 7908 4169 7936
rect 4028 7896 4034 7908
rect 4157 7905 4169 7908
rect 4203 7905 4215 7939
rect 4157 7899 4215 7905
rect 4338 7896 4344 7948
rect 4396 7936 4402 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 4396 7908 4445 7936
rect 4396 7896 4402 7908
rect 4433 7905 4445 7908
rect 4479 7936 4491 7939
rect 4706 7936 4712 7948
rect 4479 7908 4712 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 5092 7936 5120 7976
rect 5169 7973 5181 8007
rect 5215 8004 5227 8007
rect 5626 8004 5632 8016
rect 5215 7976 5632 8004
rect 5215 7973 5227 7976
rect 5169 7967 5227 7973
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 8018 8004 8024 8016
rect 5736 7976 8024 8004
rect 5350 7936 5356 7948
rect 5092 7908 5356 7936
rect 5350 7896 5356 7908
rect 5408 7936 5414 7948
rect 5736 7936 5764 7976
rect 8018 7964 8024 7976
rect 8076 7964 8082 8016
rect 5408 7908 5764 7936
rect 6089 7939 6147 7945
rect 5408 7896 5414 7908
rect 6089 7905 6101 7939
rect 6135 7936 6147 7939
rect 6730 7936 6736 7948
rect 6135 7908 6736 7936
rect 6135 7905 6147 7908
rect 6089 7899 6147 7905
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 6972 7908 7205 7936
rect 6972 7896 6978 7908
rect 7193 7905 7205 7908
rect 7239 7905 7251 7939
rect 8496 7936 8524 8035
rect 9030 7936 9036 7948
rect 8496 7908 9036 7936
rect 7193 7899 7251 7905
rect 9030 7896 9036 7908
rect 9088 7936 9094 7948
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 9088 7908 9229 7936
rect 9088 7896 9094 7908
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 9306 7896 9312 7948
rect 9364 7936 9370 7948
rect 9473 7939 9531 7945
rect 9473 7936 9485 7939
rect 9364 7908 9485 7936
rect 9364 7896 9370 7908
rect 9473 7905 9485 7908
rect 9519 7905 9531 7939
rect 9473 7899 9531 7905
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7868 5687 7871
rect 5905 7871 5963 7877
rect 5905 7868 5917 7871
rect 5675 7840 5917 7868
rect 5675 7837 5687 7840
rect 5629 7831 5687 7837
rect 5905 7837 5917 7840
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 6362 7828 6368 7880
rect 6420 7828 6426 7880
rect 6454 7828 6460 7880
rect 6512 7828 6518 7880
rect 7098 7868 7104 7880
rect 6886 7840 7104 7868
rect 3421 7803 3479 7809
rect 3421 7769 3433 7803
rect 3467 7800 3479 7803
rect 3602 7800 3608 7812
rect 3467 7772 3608 7800
rect 3467 7769 3479 7772
rect 3421 7763 3479 7769
rect 3602 7760 3608 7772
rect 3660 7760 3666 7812
rect 4062 7760 4068 7812
rect 4120 7760 4126 7812
rect 5537 7803 5595 7809
rect 5537 7769 5549 7803
rect 5583 7800 5595 7803
rect 6546 7800 6552 7812
rect 5583 7772 6552 7800
rect 5583 7769 5595 7772
rect 5537 7763 5595 7769
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 3697 7735 3755 7741
rect 3697 7701 3709 7735
rect 3743 7732 3755 7735
rect 4617 7735 4675 7741
rect 4617 7732 4629 7735
rect 3743 7704 4629 7732
rect 3743 7701 3755 7704
rect 3697 7695 3755 7701
rect 4617 7701 4629 7704
rect 4663 7701 4675 7735
rect 4617 7695 4675 7701
rect 6273 7735 6331 7741
rect 6273 7701 6285 7735
rect 6319 7732 6331 7735
rect 6886 7732 6914 7840
rect 7098 7828 7104 7840
rect 7156 7828 7162 7880
rect 8110 7760 8116 7812
rect 8168 7800 8174 7812
rect 8168 7772 9260 7800
rect 8168 7760 8174 7772
rect 6319 7704 6914 7732
rect 6319 7701 6331 7704
rect 6273 7695 6331 7701
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7101 7735 7159 7741
rect 7101 7732 7113 7735
rect 7064 7704 7113 7732
rect 7064 7692 7070 7704
rect 7101 7701 7113 7704
rect 7147 7701 7159 7735
rect 7101 7695 7159 7701
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 8570 7732 8576 7744
rect 8076 7704 8576 7732
rect 8076 7692 8082 7704
rect 8570 7692 8576 7704
rect 8628 7732 8634 7744
rect 9030 7732 9036 7744
rect 8628 7704 9036 7732
rect 8628 7692 8634 7704
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9232 7732 9260 7772
rect 10594 7732 10600 7744
rect 9232 7704 10600 7732
rect 10594 7692 10600 7704
rect 10652 7692 10658 7744
rect 552 7642 11408 7664
rect 552 7590 1755 7642
rect 1807 7590 1819 7642
rect 1871 7590 1883 7642
rect 1935 7590 1947 7642
rect 1999 7590 2011 7642
rect 2063 7590 4469 7642
rect 4521 7590 4533 7642
rect 4585 7590 4597 7642
rect 4649 7590 4661 7642
rect 4713 7590 4725 7642
rect 4777 7590 7183 7642
rect 7235 7590 7247 7642
rect 7299 7590 7311 7642
rect 7363 7590 7375 7642
rect 7427 7590 7439 7642
rect 7491 7590 9897 7642
rect 9949 7590 9961 7642
rect 10013 7590 10025 7642
rect 10077 7590 10089 7642
rect 10141 7590 10153 7642
rect 10205 7590 11408 7642
rect 552 7568 11408 7590
rect 3973 7531 4031 7537
rect 3973 7497 3985 7531
rect 4019 7528 4031 7531
rect 4062 7528 4068 7540
rect 4019 7500 4068 7528
rect 4019 7497 4031 7500
rect 3973 7491 4031 7497
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 4154 7488 4160 7540
rect 4212 7488 4218 7540
rect 6181 7531 6239 7537
rect 6181 7497 6193 7531
rect 6227 7528 6239 7531
rect 6454 7528 6460 7540
rect 6227 7500 6460 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 6546 7488 6552 7540
rect 6604 7488 6610 7540
rect 7561 7531 7619 7537
rect 7561 7497 7573 7531
rect 7607 7528 7619 7531
rect 8938 7528 8944 7540
rect 7607 7500 8944 7528
rect 7607 7497 7619 7500
rect 7561 7491 7619 7497
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 9033 7531 9091 7537
rect 9033 7497 9045 7531
rect 9079 7528 9091 7531
rect 9306 7528 9312 7540
rect 9079 7500 9312 7528
rect 9079 7497 9091 7500
rect 9033 7491 9091 7497
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 3053 7463 3111 7469
rect 3053 7429 3065 7463
rect 3099 7460 3111 7463
rect 4172 7460 4200 7488
rect 3099 7432 4200 7460
rect 6932 7432 7420 7460
rect 3099 7429 3111 7432
rect 3053 7423 3111 7429
rect 3804 7401 3832 7432
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7361 3847 7395
rect 3789 7355 3847 7361
rect 4798 7352 4804 7404
rect 4856 7352 4862 7404
rect 6362 7352 6368 7404
rect 6420 7392 6426 7404
rect 6932 7401 6960 7432
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 6420 7364 6929 7392
rect 6420 7352 6426 7364
rect 6917 7361 6929 7364
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 7006 7352 7012 7404
rect 7064 7352 7070 7404
rect 1118 7284 1124 7336
rect 1176 7324 1182 7336
rect 1673 7327 1731 7333
rect 1673 7324 1685 7327
rect 1176 7296 1685 7324
rect 1176 7284 1182 7296
rect 1673 7293 1685 7296
rect 1719 7324 1731 7327
rect 3510 7324 3516 7336
rect 1719 7296 3516 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 3510 7284 3516 7296
rect 3568 7284 3574 7336
rect 3970 7284 3976 7336
rect 4028 7284 4034 7336
rect 4617 7327 4675 7333
rect 4617 7293 4629 7327
rect 4663 7324 4675 7327
rect 4706 7324 4712 7336
rect 4663 7296 4712 7324
rect 4663 7293 4675 7296
rect 4617 7287 4675 7293
rect 4706 7284 4712 7296
rect 4764 7324 4770 7336
rect 5350 7324 5356 7336
rect 4764 7296 5356 7324
rect 4764 7284 4770 7296
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 6733 7327 6791 7333
rect 6733 7293 6745 7327
rect 6779 7293 6791 7327
rect 6733 7287 6791 7293
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7324 6883 7327
rect 7098 7324 7104 7336
rect 6871 7296 7104 7324
rect 6871 7293 6883 7296
rect 6825 7287 6883 7293
rect 1940 7259 1998 7265
rect 1940 7225 1952 7259
rect 1986 7256 1998 7259
rect 2314 7256 2320 7268
rect 1986 7228 2320 7256
rect 1986 7225 1998 7228
rect 1940 7219 1998 7225
rect 2314 7216 2320 7228
rect 2372 7216 2378 7268
rect 3988 7256 4016 7284
rect 4125 7259 4183 7265
rect 4125 7256 4137 7259
rect 3988 7228 4137 7256
rect 4125 7225 4137 7228
rect 4171 7225 4183 7259
rect 4125 7219 4183 7225
rect 4338 7216 4344 7268
rect 4396 7216 4402 7268
rect 5046 7259 5104 7265
rect 5046 7256 5058 7259
rect 4540 7228 5058 7256
rect 3237 7191 3295 7197
rect 3237 7157 3249 7191
rect 3283 7188 3295 7191
rect 3602 7188 3608 7200
rect 3283 7160 3608 7188
rect 3283 7157 3295 7160
rect 3237 7151 3295 7157
rect 3602 7148 3608 7160
rect 3660 7148 3666 7200
rect 4430 7148 4436 7200
rect 4488 7188 4494 7200
rect 4540 7197 4568 7228
rect 5046 7225 5058 7228
rect 5092 7225 5104 7259
rect 5046 7219 5104 7225
rect 4525 7191 4583 7197
rect 4525 7188 4537 7191
rect 4488 7160 4537 7188
rect 4488 7148 4494 7160
rect 4525 7157 4537 7160
rect 4571 7157 4583 7191
rect 6748 7188 6776 7287
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 7392 7265 7420 7432
rect 8386 7420 8392 7472
rect 8444 7420 8450 7472
rect 8404 7392 8432 7420
rect 7944 7364 8708 7392
rect 7469 7327 7527 7333
rect 7469 7293 7481 7327
rect 7515 7324 7527 7327
rect 7742 7324 7748 7336
rect 7515 7296 7748 7324
rect 7515 7293 7527 7296
rect 7469 7287 7527 7293
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 7944 7333 7972 7364
rect 7837 7327 7895 7333
rect 7837 7293 7849 7327
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7293 7987 7327
rect 7929 7287 7987 7293
rect 7377 7259 7435 7265
rect 7377 7225 7389 7259
rect 7423 7256 7435 7259
rect 7852 7256 7880 7287
rect 8018 7284 8024 7336
rect 8076 7284 8082 7336
rect 8205 7327 8263 7333
rect 8205 7293 8217 7327
rect 8251 7324 8263 7327
rect 8294 7324 8300 7336
rect 8251 7296 8300 7324
rect 8251 7293 8263 7296
rect 8205 7287 8263 7293
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 8389 7327 8447 7333
rect 8389 7293 8401 7327
rect 8435 7293 8447 7327
rect 8389 7287 8447 7293
rect 7423 7228 7880 7256
rect 8404 7256 8432 7287
rect 8570 7284 8576 7336
rect 8628 7284 8634 7336
rect 8680 7333 8708 7364
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 10594 7352 10600 7404
rect 10652 7352 10658 7404
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 8757 7327 8815 7333
rect 8757 7293 8769 7327
rect 8803 7324 8815 7327
rect 9140 7324 9168 7352
rect 8803 7296 9168 7324
rect 9309 7327 9367 7333
rect 8803 7293 8815 7296
rect 8757 7287 8815 7293
rect 9309 7293 9321 7327
rect 9355 7293 9367 7327
rect 9309 7287 9367 7293
rect 9125 7259 9183 7265
rect 9125 7256 9137 7259
rect 8404 7228 9137 7256
rect 7423 7225 7435 7228
rect 7377 7219 7435 7225
rect 9125 7225 9137 7228
rect 9171 7225 9183 7259
rect 9324 7256 9352 7287
rect 9398 7284 9404 7336
rect 9456 7324 9462 7336
rect 9585 7327 9643 7333
rect 9585 7324 9597 7327
rect 9456 7296 9597 7324
rect 9456 7284 9462 7296
rect 9585 7293 9597 7296
rect 9631 7293 9643 7327
rect 9585 7287 9643 7293
rect 11054 7284 11060 7336
rect 11112 7284 11118 7336
rect 10045 7259 10103 7265
rect 10045 7256 10057 7259
rect 9324 7228 10057 7256
rect 9125 7219 9183 7225
rect 10045 7225 10057 7228
rect 10091 7225 10103 7259
rect 10045 7219 10103 7225
rect 8110 7188 8116 7200
rect 6748 7160 8116 7188
rect 4525 7151 4583 7157
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 9493 7191 9551 7197
rect 9493 7188 9505 7191
rect 8260 7160 9505 7188
rect 8260 7148 8266 7160
rect 9493 7157 9505 7160
rect 9539 7157 9551 7191
rect 9493 7151 9551 7157
rect 10870 7148 10876 7200
rect 10928 7148 10934 7200
rect 552 7098 11568 7120
rect 552 7046 3112 7098
rect 3164 7046 3176 7098
rect 3228 7046 3240 7098
rect 3292 7046 3304 7098
rect 3356 7046 3368 7098
rect 3420 7046 5826 7098
rect 5878 7046 5890 7098
rect 5942 7046 5954 7098
rect 6006 7046 6018 7098
rect 6070 7046 6082 7098
rect 6134 7046 8540 7098
rect 8592 7046 8604 7098
rect 8656 7046 8668 7098
rect 8720 7046 8732 7098
rect 8784 7046 8796 7098
rect 8848 7046 11254 7098
rect 11306 7046 11318 7098
rect 11370 7046 11382 7098
rect 11434 7046 11446 7098
rect 11498 7046 11510 7098
rect 11562 7046 11568 7098
rect 552 7024 11568 7046
rect 2314 6944 2320 6996
rect 2372 6944 2378 6996
rect 3421 6987 3479 6993
rect 3421 6984 3433 6987
rect 2792 6956 3433 6984
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6848 1639 6851
rect 2314 6848 2320 6860
rect 1627 6820 2320 6848
rect 1627 6817 1639 6820
rect 1581 6811 1639 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 2406 6808 2412 6860
rect 2464 6808 2470 6860
rect 2792 6857 2820 6956
rect 3421 6953 3433 6956
rect 3467 6984 3479 6987
rect 3602 6984 3608 6996
rect 3467 6956 3608 6984
rect 3467 6953 3479 6956
rect 3421 6947 3479 6953
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 8113 6987 8171 6993
rect 8113 6984 8125 6987
rect 7800 6956 8125 6984
rect 7800 6944 7806 6956
rect 8113 6953 8125 6956
rect 8159 6984 8171 6987
rect 9122 6984 9128 6996
rect 8159 6956 9128 6984
rect 8159 6953 8171 6956
rect 8113 6947 8171 6953
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 4062 6876 4068 6928
rect 4120 6916 4126 6928
rect 5166 6916 5172 6928
rect 4120 6888 5172 6916
rect 4120 6876 4126 6888
rect 2501 6851 2559 6857
rect 2501 6817 2513 6851
rect 2547 6817 2559 6851
rect 2501 6811 2559 6817
rect 2777 6851 2835 6857
rect 2777 6817 2789 6851
rect 2823 6817 2835 6851
rect 2777 6811 2835 6817
rect 1394 6740 1400 6792
rect 1452 6780 1458 6792
rect 1765 6783 1823 6789
rect 1765 6780 1777 6783
rect 1452 6752 1777 6780
rect 1452 6740 1458 6752
rect 1765 6749 1777 6752
rect 1811 6749 1823 6783
rect 1765 6743 1823 6749
rect 1854 6740 1860 6792
rect 1912 6740 1918 6792
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 2424 6780 2452 6808
rect 2087 6752 2452 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 1302 6604 1308 6656
rect 1360 6644 1366 6656
rect 1397 6647 1455 6653
rect 1397 6644 1409 6647
rect 1360 6616 1409 6644
rect 1360 6604 1366 6616
rect 1397 6613 1409 6616
rect 1443 6613 1455 6647
rect 1397 6607 1455 6613
rect 1670 6604 1676 6656
rect 1728 6644 1734 6656
rect 1964 6644 1992 6743
rect 2516 6712 2544 6811
rect 3234 6808 3240 6860
rect 3292 6808 3298 6860
rect 3513 6851 3571 6857
rect 3513 6817 3525 6851
rect 3559 6848 3571 6851
rect 3970 6848 3976 6860
rect 3559 6820 3976 6848
rect 3559 6817 3571 6820
rect 3513 6811 3571 6817
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 3050 6780 3056 6792
rect 2731 6752 3056 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 3050 6740 3056 6752
rect 3108 6780 3114 6792
rect 3528 6780 3556 6811
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 4154 6808 4160 6860
rect 4212 6808 4218 6860
rect 4356 6857 4384 6888
rect 5166 6876 5172 6888
rect 5224 6876 5230 6928
rect 8018 6916 8024 6928
rect 7314 6888 8024 6916
rect 8018 6876 8024 6888
rect 8076 6876 8082 6928
rect 8294 6916 8300 6928
rect 8220 6888 8300 6916
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6817 4399 6851
rect 4341 6811 4399 6817
rect 4525 6851 4583 6857
rect 4525 6817 4537 6851
rect 4571 6848 4583 6851
rect 4890 6848 4896 6860
rect 4571 6820 4896 6848
rect 4571 6817 4583 6820
rect 4525 6811 4583 6817
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 7650 6808 7656 6860
rect 7708 6808 7714 6860
rect 8220 6857 8248 6888
rect 8294 6876 8300 6888
rect 8352 6876 8358 6928
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6817 8263 6851
rect 8205 6811 8263 6817
rect 3108 6752 3556 6780
rect 3108 6740 3114 6752
rect 5258 6740 5264 6792
rect 5316 6780 5322 6792
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 5316 6752 5825 6780
rect 5316 6740 5322 6752
rect 5813 6749 5825 6752
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 6546 6780 6552 6792
rect 6227 6752 6552 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 3237 6715 3295 6721
rect 3237 6712 3249 6715
rect 2516 6684 3249 6712
rect 3237 6681 3249 6684
rect 3283 6681 3295 6715
rect 3237 6675 3295 6681
rect 7098 6672 7104 6724
rect 7156 6712 7162 6724
rect 8220 6712 8248 6811
rect 9030 6808 9036 6860
rect 9088 6848 9094 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9088 6820 9689 6848
rect 9088 6808 9094 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 7156 6684 8248 6712
rect 7156 6672 7162 6684
rect 9582 6672 9588 6724
rect 9640 6712 9646 6724
rect 9692 6712 9720 6811
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 9861 6851 9919 6857
rect 9861 6848 9873 6851
rect 9824 6820 9873 6848
rect 9824 6808 9830 6820
rect 9861 6817 9873 6820
rect 9907 6817 9919 6851
rect 9861 6811 9919 6817
rect 10410 6808 10416 6860
rect 10468 6848 10474 6860
rect 10870 6848 10876 6860
rect 10468 6820 10876 6848
rect 10468 6808 10474 6820
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 10229 6715 10287 6721
rect 10229 6712 10241 6715
rect 9640 6684 10241 6712
rect 9640 6672 9646 6684
rect 10229 6681 10241 6684
rect 10275 6681 10287 6715
rect 10229 6675 10287 6681
rect 1728 6616 1992 6644
rect 1728 6604 1734 6616
rect 2222 6604 2228 6656
rect 2280 6604 2286 6656
rect 3970 6604 3976 6656
rect 4028 6604 4034 6656
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 4433 6647 4491 6653
rect 4433 6644 4445 6647
rect 4304 6616 4445 6644
rect 4304 6604 4310 6616
rect 4433 6613 4445 6616
rect 4479 6613 4491 6647
rect 4433 6607 4491 6613
rect 7837 6647 7895 6653
rect 7837 6613 7849 6647
rect 7883 6644 7895 6647
rect 8202 6644 8208 6656
rect 7883 6616 8208 6644
rect 7883 6613 7895 6616
rect 7837 6607 7895 6613
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8297 6647 8355 6653
rect 8297 6613 8309 6647
rect 8343 6644 8355 6647
rect 8386 6644 8392 6656
rect 8343 6616 8392 6644
rect 8343 6613 8355 6616
rect 8297 6607 8355 6613
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 9769 6647 9827 6653
rect 9769 6644 9781 6647
rect 9732 6616 9781 6644
rect 9732 6604 9738 6616
rect 9769 6613 9781 6616
rect 9815 6613 9827 6647
rect 9769 6607 9827 6613
rect 552 6554 11408 6576
rect 552 6502 1755 6554
rect 1807 6502 1819 6554
rect 1871 6502 1883 6554
rect 1935 6502 1947 6554
rect 1999 6502 2011 6554
rect 2063 6502 4469 6554
rect 4521 6502 4533 6554
rect 4585 6502 4597 6554
rect 4649 6502 4661 6554
rect 4713 6502 4725 6554
rect 4777 6502 7183 6554
rect 7235 6502 7247 6554
rect 7299 6502 7311 6554
rect 7363 6502 7375 6554
rect 7427 6502 7439 6554
rect 7491 6502 9897 6554
rect 9949 6502 9961 6554
rect 10013 6502 10025 6554
rect 10077 6502 10089 6554
rect 10141 6502 10153 6554
rect 10205 6502 11408 6554
rect 552 6480 11408 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 1452 6412 2176 6440
rect 1452 6400 1458 6412
rect 2148 6372 2176 6412
rect 2222 6400 2228 6452
rect 2280 6440 2286 6452
rect 2685 6443 2743 6449
rect 2685 6440 2697 6443
rect 2280 6412 2697 6440
rect 2280 6400 2286 6412
rect 2685 6409 2697 6412
rect 2731 6409 2743 6443
rect 2685 6403 2743 6409
rect 3234 6400 3240 6452
rect 3292 6440 3298 6452
rect 3878 6440 3884 6452
rect 3292 6412 3884 6440
rect 3292 6400 3298 6412
rect 3878 6400 3884 6412
rect 3936 6440 3942 6452
rect 4338 6440 4344 6452
rect 3936 6412 4344 6440
rect 3936 6400 3942 6412
rect 4338 6400 4344 6412
rect 4396 6400 4402 6452
rect 5258 6400 5264 6452
rect 5316 6400 5322 6452
rect 5350 6400 5356 6452
rect 5408 6440 5414 6452
rect 6273 6443 6331 6449
rect 6273 6440 6285 6443
rect 5408 6412 6285 6440
rect 5408 6400 5414 6412
rect 6273 6409 6285 6412
rect 6319 6440 6331 6443
rect 6822 6440 6828 6452
rect 6319 6412 6828 6440
rect 6319 6409 6331 6412
rect 6273 6403 6331 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 7650 6400 7656 6452
rect 7708 6400 7714 6452
rect 2406 6372 2412 6384
rect 2148 6344 2412 6372
rect 2406 6332 2412 6344
rect 2464 6332 2470 6384
rect 2501 6375 2559 6381
rect 2501 6341 2513 6375
rect 2547 6341 2559 6375
rect 2501 6335 2559 6341
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 2516 6304 2544 6335
rect 3050 6332 3056 6384
rect 3108 6332 3114 6384
rect 4890 6332 4896 6384
rect 4948 6372 4954 6384
rect 4948 6344 5396 6372
rect 4948 6332 4954 6344
rect 5258 6304 5264 6316
rect 2372 6276 2544 6304
rect 5092 6276 5264 6304
rect 2372 6264 2378 6276
rect 1029 6239 1087 6245
rect 1029 6205 1041 6239
rect 1075 6236 1087 6239
rect 1118 6236 1124 6248
rect 1075 6208 1124 6236
rect 1075 6205 1087 6208
rect 1029 6199 1087 6205
rect 1118 6196 1124 6208
rect 1176 6196 1182 6248
rect 1302 6245 1308 6248
rect 1296 6236 1308 6245
rect 1263 6208 1308 6236
rect 1296 6199 1308 6208
rect 1302 6196 1308 6199
rect 1360 6196 1366 6248
rect 5092 6245 5120 6276
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 5368 6304 5396 6344
rect 5368 6276 5672 6304
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6205 5135 6239
rect 5077 6199 5135 6205
rect 5166 6196 5172 6248
rect 5224 6196 5230 6248
rect 5368 6245 5396 6276
rect 5644 6245 5672 6276
rect 5353 6239 5411 6245
rect 5353 6205 5365 6239
rect 5399 6205 5411 6239
rect 5353 6199 5411 6205
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6205 5503 6239
rect 5445 6199 5503 6205
rect 5629 6239 5687 6245
rect 5629 6205 5641 6239
rect 5675 6205 5687 6239
rect 5629 6199 5687 6205
rect 3510 6128 3516 6180
rect 3568 6128 3574 6180
rect 5184 6168 5212 6196
rect 5460 6168 5488 6199
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7837 6239 7895 6245
rect 7837 6236 7849 6239
rect 6972 6208 7849 6236
rect 6972 6196 6978 6208
rect 7837 6205 7849 6208
rect 7883 6205 7895 6239
rect 7837 6199 7895 6205
rect 8113 6239 8171 6245
rect 8113 6205 8125 6239
rect 8159 6236 8171 6239
rect 8294 6236 8300 6248
rect 8159 6208 8300 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 8294 6196 8300 6208
rect 8352 6196 8358 6248
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 5184 6140 5488 6168
rect 7558 6128 7564 6180
rect 7616 6128 7622 6180
rect 8588 6168 8616 6199
rect 8938 6196 8944 6248
rect 8996 6196 9002 6248
rect 10410 6196 10416 6248
rect 10468 6196 10474 6248
rect 7760 6140 8616 6168
rect 2685 6103 2743 6109
rect 2685 6069 2697 6103
rect 2731 6100 2743 6103
rect 2866 6100 2872 6112
rect 2731 6072 2872 6100
rect 2731 6069 2743 6072
rect 2685 6063 2743 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6100 5687 6103
rect 7760 6100 7788 6140
rect 9674 6128 9680 6180
rect 9732 6128 9738 6180
rect 5675 6072 7788 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 8021 6103 8079 6109
rect 8021 6100 8033 6103
rect 7892 6072 8033 6100
rect 7892 6060 7898 6072
rect 8021 6069 8033 6072
rect 8067 6069 8079 6103
rect 8021 6063 8079 6069
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 10973 6103 11031 6109
rect 10973 6100 10985 6103
rect 9824 6072 10985 6100
rect 9824 6060 9830 6072
rect 10973 6069 10985 6072
rect 11019 6069 11031 6103
rect 10973 6063 11031 6069
rect 552 6010 11568 6032
rect 552 5958 3112 6010
rect 3164 5958 3176 6010
rect 3228 5958 3240 6010
rect 3292 5958 3304 6010
rect 3356 5958 3368 6010
rect 3420 5958 5826 6010
rect 5878 5958 5890 6010
rect 5942 5958 5954 6010
rect 6006 5958 6018 6010
rect 6070 5958 6082 6010
rect 6134 5958 8540 6010
rect 8592 5958 8604 6010
rect 8656 5958 8668 6010
rect 8720 5958 8732 6010
rect 8784 5958 8796 6010
rect 8848 5958 11254 6010
rect 11306 5958 11318 6010
rect 11370 5958 11382 6010
rect 11434 5958 11446 6010
rect 11498 5958 11510 6010
rect 11562 5958 11568 6010
rect 552 5936 11568 5958
rect 2130 5856 2136 5908
rect 2188 5896 2194 5908
rect 2501 5899 2559 5905
rect 2501 5896 2513 5899
rect 2188 5868 2513 5896
rect 2188 5856 2194 5868
rect 2501 5865 2513 5868
rect 2547 5865 2559 5899
rect 2501 5859 2559 5865
rect 2590 5856 2596 5908
rect 2648 5896 2654 5908
rect 2685 5899 2743 5905
rect 2685 5896 2697 5899
rect 2648 5868 2697 5896
rect 2648 5856 2654 5868
rect 2685 5865 2697 5868
rect 2731 5865 2743 5899
rect 2685 5859 2743 5865
rect 2869 5899 2927 5905
rect 2869 5865 2881 5899
rect 2915 5896 2927 5899
rect 2958 5896 2964 5908
rect 2915 5868 2964 5896
rect 2915 5865 2927 5868
rect 2869 5859 2927 5865
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 4890 5856 4896 5908
rect 4948 5856 4954 5908
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 5224 5868 5396 5896
rect 5224 5856 5230 5868
rect 2317 5831 2375 5837
rect 2317 5797 2329 5831
rect 2363 5828 2375 5831
rect 2406 5828 2412 5840
rect 2363 5800 2412 5828
rect 2363 5797 2375 5800
rect 2317 5791 2375 5797
rect 2406 5788 2412 5800
rect 2464 5788 2470 5840
rect 3780 5831 3838 5837
rect 3780 5797 3792 5831
rect 3826 5828 3838 5831
rect 3970 5828 3976 5840
rect 3826 5800 3976 5828
rect 3826 5797 3838 5800
rect 3780 5791 3838 5797
rect 3970 5788 3976 5800
rect 4028 5788 4034 5840
rect 1670 5720 1676 5772
rect 1728 5760 1734 5772
rect 2593 5763 2651 5769
rect 2593 5760 2605 5763
rect 1728 5732 2605 5760
rect 1728 5720 1734 5732
rect 2593 5729 2605 5732
rect 2639 5729 2651 5763
rect 2593 5723 2651 5729
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 2961 5763 3019 5769
rect 2961 5760 2973 5763
rect 2832 5732 2973 5760
rect 2832 5720 2838 5732
rect 2961 5729 2973 5732
rect 3007 5729 3019 5763
rect 4798 5760 4804 5772
rect 2961 5723 3019 5729
rect 3252 5732 4804 5760
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 1360 5664 1409 5692
rect 1360 5652 1366 5664
rect 1397 5661 1409 5664
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 2866 5652 2872 5704
rect 2924 5692 2930 5704
rect 3252 5701 3280 5732
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 4908 5760 4936 5856
rect 5368 5837 5396 5868
rect 6546 5856 6552 5908
rect 6604 5856 6610 5908
rect 7101 5899 7159 5905
rect 7101 5896 7113 5899
rect 6886 5868 7113 5896
rect 5353 5831 5411 5837
rect 5353 5797 5365 5831
rect 5399 5797 5411 5831
rect 5353 5791 5411 5797
rect 5169 5763 5227 5769
rect 5169 5760 5181 5763
rect 4908 5732 5181 5760
rect 5169 5729 5181 5732
rect 5215 5729 5227 5763
rect 5368 5758 5396 5791
rect 5445 5763 5503 5769
rect 5445 5758 5457 5763
rect 5368 5730 5457 5758
rect 5169 5723 5227 5729
rect 5445 5729 5457 5730
rect 5491 5729 5503 5763
rect 5445 5723 5503 5729
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5729 5687 5763
rect 5629 5723 5687 5729
rect 6733 5763 6791 5769
rect 6733 5729 6745 5763
rect 6779 5760 6791 5763
rect 6886 5760 6914 5868
rect 7101 5865 7113 5868
rect 7147 5865 7159 5899
rect 7101 5859 7159 5865
rect 7561 5899 7619 5905
rect 7561 5865 7573 5899
rect 7607 5896 7619 5899
rect 7742 5896 7748 5908
rect 7607 5868 7748 5896
rect 7607 5865 7619 5868
rect 7561 5859 7619 5865
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 8018 5856 8024 5908
rect 8076 5856 8082 5908
rect 8294 5856 8300 5908
rect 8352 5856 8358 5908
rect 6779 5732 6914 5760
rect 7469 5763 7527 5769
rect 6779 5729 6791 5732
rect 6733 5723 6791 5729
rect 7469 5729 7481 5763
rect 7515 5760 7527 5763
rect 7650 5760 7656 5772
rect 7515 5732 7656 5760
rect 7515 5729 7527 5732
rect 7469 5723 7527 5729
rect 3237 5695 3295 5701
rect 3237 5692 3249 5695
rect 2924 5664 3249 5692
rect 2924 5652 2930 5664
rect 3237 5661 3249 5664
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 3510 5652 3516 5704
rect 3568 5652 3574 5704
rect 5184 5692 5212 5723
rect 5644 5692 5672 5723
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7760 5760 7788 5856
rect 9858 5828 9864 5840
rect 9508 5800 9864 5828
rect 7929 5763 7987 5769
rect 7929 5760 7941 5763
rect 7760 5732 7941 5760
rect 7929 5729 7941 5732
rect 7975 5729 7987 5763
rect 7929 5723 7987 5729
rect 8113 5763 8171 5769
rect 8113 5729 8125 5763
rect 8159 5729 8171 5763
rect 8113 5723 8171 5729
rect 5184 5664 5672 5692
rect 7742 5652 7748 5704
rect 7800 5652 7806 5704
rect 7834 5652 7840 5704
rect 7892 5692 7898 5704
rect 8128 5692 8156 5723
rect 8202 5720 8208 5772
rect 8260 5720 8266 5772
rect 9508 5769 9536 5800
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5729 9551 5763
rect 9493 5723 9551 5729
rect 9508 5692 9536 5723
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 9640 5732 9689 5760
rect 9640 5720 9646 5732
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 7892 5664 9536 5692
rect 7892 5652 7898 5664
rect 3053 5627 3111 5633
rect 3053 5593 3065 5627
rect 3099 5624 3111 5627
rect 3418 5624 3424 5636
rect 3099 5596 3424 5624
rect 3099 5593 3111 5596
rect 3053 5587 3111 5593
rect 3418 5584 3424 5596
rect 3476 5584 3482 5636
rect 1578 5516 1584 5568
rect 1636 5556 1642 5568
rect 2041 5559 2099 5565
rect 2041 5556 2053 5559
rect 1636 5528 2053 5556
rect 1636 5516 1642 5528
rect 2041 5525 2053 5528
rect 2087 5525 2099 5559
rect 2041 5519 2099 5525
rect 3142 5516 3148 5568
rect 3200 5516 3206 5568
rect 4982 5516 4988 5568
rect 5040 5516 5046 5568
rect 5537 5559 5595 5565
rect 5537 5525 5549 5559
rect 5583 5556 5595 5559
rect 8478 5556 8484 5568
rect 5583 5528 8484 5556
rect 5583 5525 5595 5528
rect 5537 5519 5595 5525
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 9582 5516 9588 5568
rect 9640 5516 9646 5568
rect 552 5466 11408 5488
rect 552 5414 1755 5466
rect 1807 5414 1819 5466
rect 1871 5414 1883 5466
rect 1935 5414 1947 5466
rect 1999 5414 2011 5466
rect 2063 5414 4469 5466
rect 4521 5414 4533 5466
rect 4585 5414 4597 5466
rect 4649 5414 4661 5466
rect 4713 5414 4725 5466
rect 4777 5414 7183 5466
rect 7235 5414 7247 5466
rect 7299 5414 7311 5466
rect 7363 5414 7375 5466
rect 7427 5414 7439 5466
rect 7491 5414 9897 5466
rect 9949 5414 9961 5466
rect 10013 5414 10025 5466
rect 10077 5414 10089 5466
rect 10141 5414 10153 5466
rect 10205 5414 11408 5466
rect 552 5392 11408 5414
rect 2590 5352 2596 5364
rect 1228 5324 2596 5352
rect 1228 5157 1256 5324
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 4065 5355 4123 5361
rect 4065 5321 4077 5355
rect 4111 5352 4123 5355
rect 4154 5352 4160 5364
rect 4111 5324 4160 5352
rect 4111 5321 4123 5324
rect 4065 5315 4123 5321
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 4246 5312 4252 5364
rect 4304 5312 4310 5364
rect 8113 5355 8171 5361
rect 8113 5352 8125 5355
rect 4816 5324 8125 5352
rect 1489 5287 1547 5293
rect 1489 5253 1501 5287
rect 1535 5284 1547 5287
rect 1535 5256 2176 5284
rect 1535 5253 1547 5256
rect 1489 5247 1547 5253
rect 2148 5225 2176 5256
rect 2866 5244 2872 5296
rect 2924 5284 2930 5296
rect 3237 5287 3295 5293
rect 3237 5284 3249 5287
rect 2924 5256 3249 5284
rect 2924 5244 2930 5256
rect 3237 5253 3249 5256
rect 3283 5253 3295 5287
rect 3237 5247 3295 5253
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2222 5176 2228 5228
rect 2280 5216 2286 5228
rect 2317 5219 2375 5225
rect 2317 5216 2329 5219
rect 2280 5188 2329 5216
rect 2280 5176 2286 5188
rect 2317 5185 2329 5188
rect 2363 5185 2375 5219
rect 4264 5216 4292 5312
rect 4709 5219 4767 5225
rect 4709 5216 4721 5219
rect 4264 5188 4721 5216
rect 2317 5179 2375 5185
rect 4709 5185 4721 5188
rect 4755 5185 4767 5219
rect 4816 5216 4844 5324
rect 8113 5321 8125 5324
rect 8159 5321 8171 5355
rect 8113 5315 8171 5321
rect 9490 5312 9496 5364
rect 9548 5352 9554 5364
rect 10781 5355 10839 5361
rect 10781 5352 10793 5355
rect 9548 5324 10793 5352
rect 9548 5312 9554 5324
rect 10781 5321 10793 5324
rect 10827 5321 10839 5355
rect 10781 5315 10839 5321
rect 6362 5244 6368 5296
rect 6420 5284 6426 5296
rect 6420 5256 7604 5284
rect 6420 5244 6426 5256
rect 5077 5219 5135 5225
rect 5077 5216 5089 5219
rect 4816 5188 5089 5216
rect 4709 5179 4767 5185
rect 5077 5185 5089 5188
rect 5123 5185 5135 5219
rect 5077 5179 5135 5185
rect 1213 5151 1271 5157
rect 1213 5117 1225 5151
rect 1259 5117 1271 5151
rect 1213 5111 1271 5117
rect 1305 5151 1363 5157
rect 1305 5117 1317 5151
rect 1351 5148 1363 5151
rect 2774 5148 2780 5160
rect 1351 5120 2780 5148
rect 1351 5117 1363 5120
rect 1305 5111 1363 5117
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 3142 5108 3148 5160
rect 3200 5148 3206 5160
rect 3237 5151 3295 5157
rect 3237 5148 3249 5151
rect 3200 5120 3249 5148
rect 3200 5108 3206 5120
rect 3237 5117 3249 5120
rect 3283 5117 3295 5151
rect 3237 5111 3295 5117
rect 3418 5108 3424 5160
rect 3476 5148 3482 5160
rect 3513 5151 3571 5157
rect 3513 5148 3525 5151
rect 3476 5120 3525 5148
rect 3476 5108 3482 5120
rect 3513 5117 3525 5120
rect 3559 5148 3571 5151
rect 3602 5148 3608 5160
rect 3559 5120 3608 5148
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 3602 5108 3608 5120
rect 3660 5108 3666 5160
rect 7576 5157 7604 5256
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 7708 5188 7972 5216
rect 7708 5176 7714 5188
rect 7742 5157 7748 5160
rect 6549 5151 6607 5157
rect 6549 5117 6561 5151
rect 6595 5148 6607 5151
rect 7101 5151 7159 5157
rect 7101 5148 7113 5151
rect 6595 5120 7113 5148
rect 6595 5117 6607 5120
rect 6549 5111 6607 5117
rect 7101 5117 7113 5120
rect 7147 5117 7159 5151
rect 7101 5111 7159 5117
rect 7285 5151 7343 5157
rect 7285 5117 7297 5151
rect 7331 5117 7343 5151
rect 7285 5111 7343 5117
rect 7561 5151 7619 5157
rect 7561 5117 7573 5151
rect 7607 5117 7619 5151
rect 7740 5148 7748 5157
rect 7703 5120 7748 5148
rect 7561 5111 7619 5117
rect 7740 5111 7748 5120
rect 1489 5083 1547 5089
rect 1489 5049 1501 5083
rect 1535 5080 1547 5083
rect 2961 5083 3019 5089
rect 2961 5080 2973 5083
rect 1535 5052 2973 5080
rect 1535 5049 1547 5052
rect 1489 5043 1547 5049
rect 2961 5049 2973 5052
rect 3007 5080 3019 5083
rect 3878 5080 3884 5092
rect 3007 5052 3884 5080
rect 3007 5049 3019 5052
rect 2961 5043 3019 5049
rect 3878 5040 3884 5052
rect 3936 5040 3942 5092
rect 4433 5083 4491 5089
rect 4433 5049 4445 5083
rect 4479 5080 4491 5083
rect 4706 5080 4712 5092
rect 4479 5052 4712 5080
rect 4479 5049 4491 5052
rect 4433 5043 4491 5049
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 6178 5040 6184 5092
rect 6236 5040 6242 5092
rect 6914 5040 6920 5092
rect 6972 5080 6978 5092
rect 7300 5080 7328 5111
rect 7742 5108 7748 5111
rect 7800 5108 7806 5160
rect 7944 5157 7972 5188
rect 8478 5176 8484 5228
rect 8536 5176 8542 5228
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5117 7987 5151
rect 8294 5148 8300 5160
rect 7929 5111 7987 5117
rect 8036 5120 8300 5148
rect 6972 5052 7328 5080
rect 7837 5083 7895 5089
rect 6972 5040 6978 5052
rect 7837 5049 7849 5083
rect 7883 5080 7895 5083
rect 8036 5080 8064 5120
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 8386 5108 8392 5160
rect 8444 5148 8450 5160
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 8444 5120 8861 5148
rect 8444 5108 8450 5120
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 10321 5151 10379 5157
rect 10321 5117 10333 5151
rect 10367 5148 10379 5151
rect 10410 5148 10416 5160
rect 10367 5120 10416 5148
rect 10367 5117 10379 5120
rect 10321 5111 10379 5117
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 7883 5052 8064 5080
rect 7883 5049 7895 5052
rect 7837 5043 7895 5049
rect 8110 5040 8116 5092
rect 8168 5040 8174 5092
rect 9582 5040 9588 5092
rect 9640 5040 9646 5092
rect 1394 4972 1400 5024
rect 1452 5012 1458 5024
rect 1581 5015 1639 5021
rect 1581 5012 1593 5015
rect 1452 4984 1593 5012
rect 1452 4972 1458 4984
rect 1581 4981 1593 4984
rect 1627 4981 1639 5015
rect 1581 4975 1639 4981
rect 2774 4972 2780 5024
rect 2832 5012 2838 5024
rect 3421 5015 3479 5021
rect 3421 5012 3433 5015
rect 2832 4984 3433 5012
rect 2832 4972 2838 4984
rect 3421 4981 3433 4984
rect 3467 4981 3479 5015
rect 3421 4975 3479 4981
rect 4233 5015 4291 5021
rect 4233 4981 4245 5015
rect 4279 5012 4291 5015
rect 4982 5012 4988 5024
rect 4279 4984 4988 5012
rect 4279 4981 4291 4984
rect 4233 4975 4291 4981
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 6733 5015 6791 5021
rect 6733 4981 6745 5015
rect 6779 5012 6791 5015
rect 6822 5012 6828 5024
rect 6779 4984 6828 5012
rect 6779 4981 6791 4984
rect 6733 4975 6791 4981
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 7006 4972 7012 5024
rect 7064 4972 7070 5024
rect 7466 4972 7472 5024
rect 7524 4972 7530 5024
rect 10226 4972 10232 5024
rect 10284 5012 10290 5024
rect 10505 5015 10563 5021
rect 10505 5012 10517 5015
rect 10284 4984 10517 5012
rect 10284 4972 10290 4984
rect 10505 4981 10517 4984
rect 10551 4981 10563 5015
rect 10505 4975 10563 4981
rect 552 4922 11568 4944
rect 552 4870 3112 4922
rect 3164 4870 3176 4922
rect 3228 4870 3240 4922
rect 3292 4870 3304 4922
rect 3356 4870 3368 4922
rect 3420 4870 5826 4922
rect 5878 4870 5890 4922
rect 5942 4870 5954 4922
rect 6006 4870 6018 4922
rect 6070 4870 6082 4922
rect 6134 4870 8540 4922
rect 8592 4870 8604 4922
rect 8656 4870 8668 4922
rect 8720 4870 8732 4922
rect 8784 4870 8796 4922
rect 8848 4870 11254 4922
rect 11306 4870 11318 4922
rect 11370 4870 11382 4922
rect 11434 4870 11446 4922
rect 11498 4870 11510 4922
rect 11562 4870 11568 4922
rect 552 4848 11568 4870
rect 1121 4811 1179 4817
rect 1121 4777 1133 4811
rect 1167 4808 1179 4811
rect 1302 4808 1308 4820
rect 1167 4780 1308 4808
rect 1167 4777 1179 4780
rect 1121 4771 1179 4777
rect 1302 4768 1308 4780
rect 1360 4768 1366 4820
rect 2222 4768 2228 4820
rect 2280 4808 2286 4820
rect 2685 4811 2743 4817
rect 2685 4808 2697 4811
rect 2280 4780 2697 4808
rect 2280 4768 2286 4780
rect 2685 4777 2697 4780
rect 2731 4777 2743 4811
rect 2685 4771 2743 4777
rect 2774 4768 2780 4820
rect 2832 4768 2838 4820
rect 6178 4768 6184 4820
rect 6236 4808 6242 4820
rect 6273 4811 6331 4817
rect 6273 4808 6285 4811
rect 6236 4780 6285 4808
rect 6236 4768 6242 4780
rect 6273 4777 6285 4780
rect 6319 4777 6331 4811
rect 6273 4771 6331 4777
rect 6917 4811 6975 4817
rect 6917 4777 6929 4811
rect 6963 4808 6975 4811
rect 7466 4808 7472 4820
rect 6963 4780 7472 4808
rect 6963 4777 6975 4780
rect 6917 4771 6975 4777
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 8110 4768 8116 4820
rect 8168 4808 8174 4820
rect 8481 4811 8539 4817
rect 8481 4808 8493 4811
rect 8168 4780 8493 4808
rect 8168 4768 8174 4780
rect 8481 4777 8493 4780
rect 8527 4777 8539 4811
rect 8481 4771 8539 4777
rect 1394 4740 1400 4752
rect 1044 4712 1400 4740
rect 1044 4681 1072 4712
rect 1394 4700 1400 4712
rect 1452 4700 1458 4752
rect 1578 4749 1584 4752
rect 1572 4740 1584 4749
rect 1539 4712 1584 4740
rect 1572 4703 1584 4712
rect 1578 4700 1584 4703
rect 1636 4700 1642 4752
rect 2590 4700 2596 4752
rect 2648 4740 2654 4752
rect 3786 4740 3792 4752
rect 2648 4712 3792 4740
rect 2648 4700 2654 4712
rect 3712 4681 3740 4712
rect 3786 4700 3792 4712
rect 3844 4700 3850 4752
rect 7006 4740 7012 4752
rect 6288 4712 7012 4740
rect 1029 4675 1087 4681
rect 1029 4641 1041 4675
rect 1075 4641 1087 4675
rect 1029 4635 1087 4641
rect 1213 4675 1271 4681
rect 1213 4641 1225 4675
rect 1259 4672 1271 4675
rect 3697 4675 3755 4681
rect 1259 4644 3556 4672
rect 1259 4641 1271 4644
rect 1213 4635 1271 4641
rect 1118 4564 1124 4616
rect 1176 4604 1182 4616
rect 3528 4613 3556 4644
rect 3697 4641 3709 4675
rect 3743 4641 3755 4675
rect 3697 4635 3755 4641
rect 3878 4632 3884 4684
rect 3936 4632 3942 4684
rect 6288 4681 6316 4712
rect 7006 4700 7012 4712
rect 7064 4700 7070 4752
rect 8849 4743 8907 4749
rect 8849 4709 8861 4743
rect 8895 4740 8907 4743
rect 10226 4740 10232 4752
rect 8895 4712 10232 4740
rect 8895 4709 8907 4712
rect 8849 4703 8907 4709
rect 10226 4700 10232 4712
rect 10284 4700 10290 4752
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4641 6331 4675
rect 6273 4635 6331 4641
rect 6362 4632 6368 4684
rect 6420 4672 6426 4684
rect 6457 4675 6515 4681
rect 6457 4672 6469 4675
rect 6420 4644 6469 4672
rect 6420 4632 6426 4644
rect 6457 4641 6469 4644
rect 6503 4641 6515 4675
rect 6457 4635 6515 4641
rect 6822 4632 6828 4684
rect 6880 4632 6886 4684
rect 8941 4675 8999 4681
rect 8941 4641 8953 4675
rect 8987 4672 8999 4675
rect 9122 4672 9128 4684
rect 8987 4644 9128 4672
rect 8987 4641 8999 4644
rect 8941 4635 8999 4641
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 1305 4607 1363 4613
rect 1305 4604 1317 4607
rect 1176 4576 1317 4604
rect 1176 4564 1182 4576
rect 1305 4573 1317 4576
rect 1351 4573 1363 4607
rect 3329 4607 3387 4613
rect 3329 4604 3341 4607
rect 1305 4567 1363 4573
rect 2700 4576 3341 4604
rect 1670 4428 1676 4480
rect 1728 4468 1734 4480
rect 2700 4468 2728 4576
rect 3329 4573 3341 4576
rect 3375 4573 3387 4607
rect 3329 4567 3387 4573
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 3344 4536 3372 4567
rect 3804 4536 3832 4567
rect 3970 4564 3976 4616
rect 4028 4564 4034 4616
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4604 9091 4607
rect 9674 4604 9680 4616
rect 9079 4576 9680 4604
rect 9079 4573 9091 4576
rect 9033 4567 9091 4573
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 3344 4508 3832 4536
rect 1728 4440 2728 4468
rect 1728 4428 1734 4440
rect 552 4378 11408 4400
rect 552 4326 1755 4378
rect 1807 4326 1819 4378
rect 1871 4326 1883 4378
rect 1935 4326 1947 4378
rect 1999 4326 2011 4378
rect 2063 4326 4469 4378
rect 4521 4326 4533 4378
rect 4585 4326 4597 4378
rect 4649 4326 4661 4378
rect 4713 4326 4725 4378
rect 4777 4326 7183 4378
rect 7235 4326 7247 4378
rect 7299 4326 7311 4378
rect 7363 4326 7375 4378
rect 7427 4326 7439 4378
rect 7491 4326 9897 4378
rect 9949 4326 9961 4378
rect 10013 4326 10025 4378
rect 10077 4326 10089 4378
rect 10141 4326 10153 4378
rect 10205 4326 11408 4378
rect 552 4304 11408 4326
rect 1670 4224 1676 4276
rect 1728 4224 1734 4276
rect 7101 4267 7159 4273
rect 7101 4233 7113 4267
rect 7147 4264 7159 4267
rect 7742 4264 7748 4276
rect 7147 4236 7748 4264
rect 7147 4233 7159 4236
rect 7101 4227 7159 4233
rect 7742 4224 7748 4236
rect 7800 4224 7806 4276
rect 9766 4224 9772 4276
rect 9824 4224 9830 4276
rect 7650 4156 7656 4208
rect 7708 4156 7714 4208
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 4028 4100 5672 4128
rect 4028 4088 4034 4100
rect 5644 4072 5672 4100
rect 7300 4100 8248 4128
rect 2786 4063 2844 4069
rect 2786 4029 2798 4063
rect 2832 4029 2844 4063
rect 2786 4023 2844 4029
rect 2792 3992 2820 4023
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 3053 4063 3111 4069
rect 3053 4060 3065 4063
rect 3016 4032 3065 4060
rect 3016 4020 3022 4032
rect 3053 4029 3065 4032
rect 3099 4060 3111 4063
rect 3510 4060 3516 4072
rect 3099 4032 3516 4060
rect 3099 4029 3111 4032
rect 3053 4023 3111 4029
rect 3510 4020 3516 4032
rect 3568 4020 3574 4072
rect 4246 4020 4252 4072
rect 4304 4060 4310 4072
rect 4709 4063 4767 4069
rect 4709 4060 4721 4063
rect 4304 4032 4721 4060
rect 4304 4020 4310 4032
rect 4709 4029 4721 4032
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 5626 4020 5632 4072
rect 5684 4060 5690 4072
rect 5905 4063 5963 4069
rect 5905 4060 5917 4063
rect 5684 4032 5917 4060
rect 5684 4020 5690 4032
rect 5905 4029 5917 4032
rect 5951 4029 5963 4063
rect 5905 4023 5963 4029
rect 6089 4063 6147 4069
rect 6089 4029 6101 4063
rect 6135 4060 6147 4063
rect 6362 4060 6368 4072
rect 6135 4032 6368 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 6362 4020 6368 4032
rect 6420 4020 6426 4072
rect 7300 4069 7328 4100
rect 8220 4072 8248 4100
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 8352 4100 8401 4128
rect 8352 4088 8358 4100
rect 8389 4097 8401 4100
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 8996 4100 9505 4128
rect 8996 4088 9002 4100
rect 9493 4097 9505 4100
rect 9539 4097 9551 4131
rect 9493 4091 9551 4097
rect 9582 4088 9588 4140
rect 9640 4088 9646 4140
rect 7285 4063 7343 4069
rect 7285 4029 7297 4063
rect 7331 4029 7343 4063
rect 7285 4023 7343 4029
rect 7561 4063 7619 4069
rect 7561 4029 7573 4063
rect 7607 4060 7619 4063
rect 7742 4060 7748 4072
rect 7607 4032 7748 4060
rect 7607 4029 7619 4032
rect 7561 4023 7619 4029
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 7837 4063 7895 4069
rect 7837 4029 7849 4063
rect 7883 4060 7895 4063
rect 7926 4060 7932 4072
rect 7883 4032 7932 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 2866 3992 2872 4004
rect 2792 3964 2872 3992
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 7469 3995 7527 4001
rect 7469 3961 7481 3995
rect 7515 3992 7527 3995
rect 7852 3992 7880 4023
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8110 4020 8116 4072
rect 8168 4020 8174 4072
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 8573 4063 8631 4069
rect 8573 4060 8585 4063
rect 8260 4032 8585 4060
rect 8260 4020 8266 4032
rect 8573 4029 8585 4032
rect 8619 4029 8631 4063
rect 8573 4023 8631 4029
rect 8665 4063 8723 4069
rect 8665 4029 8677 4063
rect 8711 4060 8723 4063
rect 8754 4060 8760 4072
rect 8711 4032 8760 4060
rect 8711 4029 8723 4032
rect 8665 4023 8723 4029
rect 8754 4020 8760 4032
rect 8812 4020 8818 4072
rect 8849 4063 8907 4069
rect 8849 4029 8861 4063
rect 8895 4029 8907 4063
rect 8849 4023 8907 4029
rect 7515 3964 7880 3992
rect 8389 3995 8447 4001
rect 7515 3961 7527 3964
rect 7469 3955 7527 3961
rect 8389 3961 8401 3995
rect 8435 3992 8447 3995
rect 8864 3992 8892 4023
rect 9030 4020 9036 4072
rect 9088 4020 9094 4072
rect 9122 4020 9128 4072
rect 9180 4020 9186 4072
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4060 9275 4063
rect 9306 4060 9312 4072
rect 9263 4032 9312 4060
rect 9263 4029 9275 4032
rect 9217 4023 9275 4029
rect 9306 4020 9312 4032
rect 9364 4060 9370 4072
rect 9766 4060 9772 4072
rect 9364 4032 9772 4060
rect 9364 4020 9370 4032
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4029 9919 4063
rect 9861 4023 9919 4029
rect 8435 3964 8892 3992
rect 9140 3992 9168 4020
rect 9585 3995 9643 4001
rect 9585 3992 9597 3995
rect 9140 3964 9597 3992
rect 8435 3961 8447 3964
rect 8389 3955 8447 3961
rect 9585 3961 9597 3964
rect 9631 3961 9643 3995
rect 9876 3992 9904 4023
rect 9585 3955 9643 3961
rect 9784 3964 9904 3992
rect 4798 3884 4804 3936
rect 4856 3884 4862 3936
rect 5997 3927 6055 3933
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 6178 3924 6184 3936
rect 6043 3896 6184 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 6178 3884 6184 3896
rect 6236 3924 6242 3936
rect 6914 3924 6920 3936
rect 6236 3896 6920 3924
rect 6236 3884 6242 3896
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 8018 3884 8024 3936
rect 8076 3924 8082 3936
rect 9784 3924 9812 3964
rect 8076 3896 9812 3924
rect 8076 3884 8082 3896
rect 552 3834 11568 3856
rect 552 3782 3112 3834
rect 3164 3782 3176 3834
rect 3228 3782 3240 3834
rect 3292 3782 3304 3834
rect 3356 3782 3368 3834
rect 3420 3782 5826 3834
rect 5878 3782 5890 3834
rect 5942 3782 5954 3834
rect 6006 3782 6018 3834
rect 6070 3782 6082 3834
rect 6134 3782 8540 3834
rect 8592 3782 8604 3834
rect 8656 3782 8668 3834
rect 8720 3782 8732 3834
rect 8784 3782 8796 3834
rect 8848 3782 11254 3834
rect 11306 3782 11318 3834
rect 11370 3782 11382 3834
rect 11434 3782 11446 3834
rect 11498 3782 11510 3834
rect 11562 3782 11568 3834
rect 552 3760 11568 3782
rect 3697 3723 3755 3729
rect 3697 3689 3709 3723
rect 3743 3720 3755 3723
rect 3786 3720 3792 3732
rect 3743 3692 3792 3720
rect 3743 3689 3755 3692
rect 3697 3683 3755 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 8110 3680 8116 3732
rect 8168 3720 8174 3732
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 8168 3692 8493 3720
rect 8168 3680 8174 3692
rect 8481 3689 8493 3692
rect 8527 3689 8539 3723
rect 8481 3683 8539 3689
rect 9030 3680 9036 3732
rect 9088 3720 9094 3732
rect 9125 3723 9183 3729
rect 9125 3720 9137 3723
rect 9088 3692 9137 3720
rect 9088 3680 9094 3692
rect 9125 3689 9137 3692
rect 9171 3689 9183 3723
rect 9125 3683 9183 3689
rect 2958 3652 2964 3664
rect 2332 3624 2964 3652
rect 2332 3593 2360 3624
rect 2958 3612 2964 3624
rect 3016 3612 3022 3664
rect 6365 3655 6423 3661
rect 6365 3652 6377 3655
rect 6012 3624 6377 3652
rect 2590 3593 2596 3596
rect 2317 3587 2375 3593
rect 2317 3553 2329 3587
rect 2363 3553 2375 3587
rect 2317 3547 2375 3553
rect 2584 3547 2596 3593
rect 2590 3544 2596 3547
rect 2648 3544 2654 3596
rect 5718 3544 5724 3596
rect 5776 3584 5782 3596
rect 6012 3593 6040 3624
rect 6365 3621 6377 3624
rect 6411 3621 6423 3655
rect 6365 3615 6423 3621
rect 6886 3624 8156 3652
rect 5997 3587 6055 3593
rect 5997 3584 6009 3587
rect 5776 3556 6009 3584
rect 5776 3544 5782 3556
rect 5997 3553 6009 3556
rect 6043 3553 6055 3587
rect 5997 3547 6055 3553
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3584 6331 3587
rect 6638 3584 6644 3596
rect 6319 3556 6644 3584
rect 6319 3553 6331 3556
rect 6273 3547 6331 3553
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 6886 3584 6914 3624
rect 6748 3556 6914 3584
rect 6365 3519 6423 3525
rect 6365 3485 6377 3519
rect 6411 3485 6423 3519
rect 6365 3479 6423 3485
rect 6181 3451 6239 3457
rect 6181 3417 6193 3451
rect 6227 3448 6239 3451
rect 6380 3448 6408 3479
rect 6227 3420 6408 3448
rect 6227 3417 6239 3420
rect 6181 3411 6239 3417
rect 4890 3340 4896 3392
rect 4948 3380 4954 3392
rect 5813 3383 5871 3389
rect 5813 3380 5825 3383
rect 4948 3352 5825 3380
rect 4948 3340 4954 3352
rect 5813 3349 5825 3352
rect 5859 3349 5871 3383
rect 6380 3380 6408 3420
rect 6549 3451 6607 3457
rect 6549 3417 6561 3451
rect 6595 3448 6607 3451
rect 6748 3448 6776 3556
rect 7742 3544 7748 3596
rect 7800 3544 7806 3596
rect 7926 3544 7932 3596
rect 7984 3544 7990 3596
rect 8128 3593 8156 3624
rect 8386 3612 8392 3664
rect 8444 3612 8450 3664
rect 8680 3624 10272 3652
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3584 8171 3587
rect 8202 3584 8208 3596
rect 8159 3556 8208 3584
rect 8159 3553 8171 3556
rect 8113 3547 8171 3553
rect 8202 3544 8208 3556
rect 8260 3584 8266 3596
rect 8478 3584 8484 3596
rect 8260 3556 8484 3584
rect 8260 3544 8266 3556
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 8680 3593 8708 3624
rect 10244 3596 10272 3624
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3553 8723 3587
rect 8665 3547 8723 3553
rect 8941 3587 8999 3593
rect 8941 3553 8953 3587
rect 8987 3584 8999 3587
rect 9030 3584 9036 3596
rect 8987 3556 9036 3584
rect 8987 3553 8999 3556
rect 8941 3547 8999 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 9306 3544 9312 3596
rect 9364 3544 9370 3596
rect 9493 3587 9551 3593
rect 9493 3553 9505 3587
rect 9539 3553 9551 3587
rect 9493 3547 9551 3553
rect 7837 3519 7895 3525
rect 7837 3516 7849 3519
rect 6886 3508 7849 3516
rect 6595 3420 6776 3448
rect 6840 3488 7849 3508
rect 6840 3480 6914 3488
rect 7837 3485 7849 3488
rect 7883 3516 7895 3519
rect 8294 3516 8300 3528
rect 7883 3488 8300 3516
rect 7883 3485 7895 3488
rect 6595 3417 6607 3420
rect 6549 3411 6607 3417
rect 6840 3380 6868 3480
rect 7837 3479 7895 3485
rect 8294 3476 8300 3488
rect 8352 3516 8358 3528
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 8352 3488 8401 3516
rect 8352 3476 8358 3488
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8570 3476 8576 3528
rect 8628 3516 8634 3528
rect 8757 3519 8815 3525
rect 8757 3516 8769 3519
rect 8628 3488 8769 3516
rect 8628 3476 8634 3488
rect 8757 3485 8769 3488
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 8849 3519 8907 3525
rect 8849 3485 8861 3519
rect 8895 3516 8907 3519
rect 9122 3516 9128 3528
rect 8895 3488 9128 3516
rect 8895 3485 8907 3488
rect 8849 3479 8907 3485
rect 9122 3476 9128 3488
rect 9180 3516 9186 3528
rect 9508 3516 9536 3547
rect 9582 3544 9588 3596
rect 9640 3544 9646 3596
rect 10226 3544 10232 3596
rect 10284 3544 10290 3596
rect 9180 3488 9536 3516
rect 10321 3519 10379 3525
rect 9180 3476 9186 3488
rect 10321 3485 10333 3519
rect 10367 3516 10379 3519
rect 10410 3516 10416 3528
rect 10367 3488 10416 3516
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 10410 3476 10416 3488
rect 10468 3476 10474 3528
rect 8205 3451 8263 3457
rect 8205 3417 8217 3451
rect 8251 3448 8263 3451
rect 9861 3451 9919 3457
rect 9861 3448 9873 3451
rect 8251 3420 9873 3448
rect 8251 3417 8263 3420
rect 8205 3411 8263 3417
rect 9861 3417 9873 3420
rect 9907 3417 9919 3451
rect 9861 3411 9919 3417
rect 6380 3352 6868 3380
rect 5813 3343 5871 3349
rect 7926 3340 7932 3392
rect 7984 3380 7990 3392
rect 9398 3380 9404 3392
rect 7984 3352 9404 3380
rect 7984 3340 7990 3352
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 552 3290 11408 3312
rect 552 3238 1755 3290
rect 1807 3238 1819 3290
rect 1871 3238 1883 3290
rect 1935 3238 1947 3290
rect 1999 3238 2011 3290
rect 2063 3238 4469 3290
rect 4521 3238 4533 3290
rect 4585 3238 4597 3290
rect 4649 3238 4661 3290
rect 4713 3238 4725 3290
rect 4777 3238 7183 3290
rect 7235 3238 7247 3290
rect 7299 3238 7311 3290
rect 7363 3238 7375 3290
rect 7427 3238 7439 3290
rect 7491 3238 9897 3290
rect 9949 3238 9961 3290
rect 10013 3238 10025 3290
rect 10077 3238 10089 3290
rect 10141 3238 10153 3290
rect 10205 3238 11408 3290
rect 552 3216 11408 3238
rect 2590 3136 2596 3188
rect 2648 3176 2654 3188
rect 2685 3179 2743 3185
rect 2685 3176 2697 3179
rect 2648 3148 2697 3176
rect 2648 3136 2654 3148
rect 2685 3145 2697 3148
rect 2731 3145 2743 3179
rect 2685 3139 2743 3145
rect 3237 3179 3295 3185
rect 3237 3145 3249 3179
rect 3283 3176 3295 3179
rect 3602 3176 3608 3188
rect 3283 3148 3608 3176
rect 3283 3145 3295 3148
rect 3237 3139 3295 3145
rect 2685 2975 2743 2981
rect 2685 2941 2697 2975
rect 2731 2941 2743 2975
rect 2685 2935 2743 2941
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 3252 2972 3280 3139
rect 3602 3136 3608 3148
rect 3660 3136 3666 3188
rect 7742 3136 7748 3188
rect 7800 3176 7806 3188
rect 8389 3179 8447 3185
rect 8389 3176 8401 3179
rect 7800 3148 8401 3176
rect 7800 3136 7806 3148
rect 8389 3145 8401 3148
rect 8435 3145 8447 3179
rect 8389 3139 8447 3145
rect 8478 3136 8484 3188
rect 8536 3176 8542 3188
rect 9033 3179 9091 3185
rect 9033 3176 9045 3179
rect 8536 3148 9045 3176
rect 8536 3136 8542 3148
rect 9033 3145 9045 3148
rect 9079 3145 9091 3179
rect 9033 3139 9091 3145
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 9456 3148 9628 3176
rect 9456 3136 9462 3148
rect 8202 3068 8208 3120
rect 8260 3108 8266 3120
rect 8846 3108 8852 3120
rect 8260 3080 8852 3108
rect 8260 3068 8266 3080
rect 8846 3068 8852 3080
rect 8904 3108 8910 3120
rect 9490 3108 9496 3120
rect 8904 3080 9496 3108
rect 8904 3068 8910 3080
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 9600 3117 9628 3148
rect 9674 3136 9680 3188
rect 9732 3136 9738 3188
rect 9858 3136 9864 3188
rect 9916 3136 9922 3188
rect 10410 3136 10416 3188
rect 10468 3136 10474 3188
rect 9585 3111 9643 3117
rect 9585 3077 9597 3111
rect 9631 3077 9643 3111
rect 9585 3071 9643 3077
rect 3786 3000 3792 3052
rect 3844 3000 3850 3052
rect 4890 3000 4896 3052
rect 4948 3000 4954 3052
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 8478 3040 8484 3052
rect 8159 3012 8484 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 2915 2944 3280 2972
rect 4617 2975 4675 2981
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 4617 2941 4629 2975
rect 4663 2941 4675 2975
rect 6178 2972 6184 2984
rect 6026 2944 6184 2972
rect 4617 2935 4675 2941
rect 2700 2904 2728 2935
rect 3970 2904 3976 2916
rect 2700 2876 3976 2904
rect 3970 2864 3976 2876
rect 4028 2864 4034 2916
rect 4632 2904 4660 2935
rect 6178 2932 6184 2944
rect 6236 2932 6242 2984
rect 6380 2972 6408 3003
rect 8478 3000 8484 3012
rect 8536 3000 8542 3052
rect 8665 3043 8723 3049
rect 8665 3009 8677 3043
rect 8711 3040 8723 3043
rect 9122 3040 9128 3052
rect 8711 3012 9128 3040
rect 8711 3009 8723 3012
rect 8665 3003 8723 3009
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 9232 3012 10272 3040
rect 6638 2972 6644 2984
rect 6380 2944 6644 2972
rect 6638 2932 6644 2944
rect 6696 2972 6702 2984
rect 8021 2975 8079 2981
rect 8021 2972 8033 2975
rect 6696 2944 8033 2972
rect 6696 2932 6702 2944
rect 8021 2941 8033 2944
rect 8067 2972 8079 2975
rect 8386 2972 8392 2984
rect 8067 2944 8392 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8386 2932 8392 2944
rect 8444 2972 8450 2984
rect 8573 2975 8631 2981
rect 8573 2972 8585 2975
rect 8444 2944 8585 2972
rect 8444 2932 8450 2944
rect 8573 2941 8585 2944
rect 8619 2941 8631 2975
rect 8757 2975 8815 2981
rect 8757 2972 8769 2975
rect 8573 2935 8631 2941
rect 8680 2944 8769 2972
rect 4798 2904 4804 2916
rect 4632 2876 4804 2904
rect 4798 2864 4804 2876
rect 4856 2864 4862 2916
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 8680 2904 8708 2944
rect 8757 2941 8769 2944
rect 8803 2941 8815 2975
rect 8757 2935 8815 2941
rect 8846 2932 8852 2984
rect 8904 2932 8910 2984
rect 9030 2932 9036 2984
rect 9088 2972 9094 2984
rect 9232 2981 9260 3012
rect 10244 2981 10272 3012
rect 9217 2975 9275 2981
rect 9217 2972 9229 2975
rect 9088 2944 9229 2972
rect 9088 2932 9094 2944
rect 9217 2941 9229 2944
rect 9263 2941 9275 2975
rect 9861 2975 9919 2981
rect 9508 2972 9628 2974
rect 9861 2972 9873 2975
rect 9217 2935 9275 2941
rect 9416 2946 9873 2972
rect 9416 2944 9536 2946
rect 9600 2944 9873 2946
rect 9309 2907 9367 2913
rect 9309 2904 9321 2907
rect 8352 2876 8708 2904
rect 8772 2876 9321 2904
rect 8352 2864 8358 2876
rect 8772 2848 8800 2876
rect 9309 2873 9321 2876
rect 9355 2873 9367 2907
rect 9309 2867 9367 2873
rect 9416 2848 9444 2944
rect 9861 2941 9873 2944
rect 9907 2941 9919 2975
rect 9861 2935 9919 2941
rect 10229 2975 10287 2981
rect 10229 2941 10241 2975
rect 10275 2941 10287 2975
rect 10229 2935 10287 2941
rect 10321 2975 10379 2981
rect 10321 2941 10333 2975
rect 10367 2941 10379 2975
rect 10505 2975 10563 2981
rect 10505 2972 10517 2975
rect 10321 2935 10379 2941
rect 10428 2944 10517 2972
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 10336 2904 10364 2935
rect 9732 2876 10364 2904
rect 9732 2864 9738 2876
rect 8754 2796 8760 2848
rect 8812 2796 8818 2848
rect 9122 2796 9128 2848
rect 9180 2836 9186 2848
rect 9398 2836 9404 2848
rect 9180 2808 9404 2836
rect 9180 2796 9186 2808
rect 9398 2796 9404 2808
rect 9456 2796 9462 2848
rect 9490 2796 9496 2848
rect 9548 2836 9554 2848
rect 10428 2836 10456 2944
rect 10505 2941 10517 2944
rect 10551 2941 10563 2975
rect 10505 2935 10563 2941
rect 9548 2808 10456 2836
rect 9548 2796 9554 2808
rect 552 2746 11568 2768
rect 552 2694 3112 2746
rect 3164 2694 3176 2746
rect 3228 2694 3240 2746
rect 3292 2694 3304 2746
rect 3356 2694 3368 2746
rect 3420 2694 5826 2746
rect 5878 2694 5890 2746
rect 5942 2694 5954 2746
rect 6006 2694 6018 2746
rect 6070 2694 6082 2746
rect 6134 2694 8540 2746
rect 8592 2694 8604 2746
rect 8656 2694 8668 2746
rect 8720 2694 8732 2746
rect 8784 2694 8796 2746
rect 8848 2694 11254 2746
rect 11306 2694 11318 2746
rect 11370 2694 11382 2746
rect 11434 2694 11446 2746
rect 11498 2694 11510 2746
rect 11562 2694 11568 2746
rect 552 2672 11568 2694
rect 6362 2592 6368 2644
rect 6420 2632 6426 2644
rect 7742 2632 7748 2644
rect 6420 2604 7748 2632
rect 6420 2592 6426 2604
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 9030 2592 9036 2644
rect 9088 2592 9094 2644
rect 9858 2632 9864 2644
rect 9416 2604 9864 2632
rect 5074 2456 5080 2508
rect 5132 2456 5138 2508
rect 5626 2456 5632 2508
rect 5684 2496 5690 2508
rect 5994 2496 6000 2508
rect 5684 2468 6000 2496
rect 5684 2456 5690 2468
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6181 2499 6239 2505
rect 6181 2465 6193 2499
rect 6227 2496 6239 2499
rect 6380 2496 6408 2592
rect 8294 2524 8300 2576
rect 8352 2524 8358 2576
rect 8386 2524 8392 2576
rect 8444 2564 8450 2576
rect 9277 2567 9335 2573
rect 9277 2564 9289 2567
rect 8444 2536 9289 2564
rect 8444 2524 8450 2536
rect 9277 2533 9289 2536
rect 9323 2564 9335 2567
rect 9416 2564 9444 2604
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 9323 2536 9444 2564
rect 9493 2567 9551 2573
rect 9323 2533 9335 2536
rect 9277 2527 9335 2533
rect 9493 2533 9505 2567
rect 9539 2533 9551 2567
rect 9493 2527 9551 2533
rect 6227 2468 6408 2496
rect 8312 2496 8340 2524
rect 9122 2496 9128 2508
rect 8312 2468 9128 2496
rect 6227 2465 6239 2468
rect 6181 2459 6239 2465
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2428 5227 2431
rect 5718 2428 5724 2440
rect 5215 2400 5724 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 8294 2388 8300 2440
rect 8352 2428 8358 2440
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 8352 2400 8585 2428
rect 8352 2388 8358 2400
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 8956 2369 8984 2468
rect 9122 2456 9128 2468
rect 9180 2496 9186 2508
rect 9508 2496 9536 2527
rect 9180 2468 9536 2496
rect 9180 2456 9186 2468
rect 8941 2363 8999 2369
rect 8941 2329 8953 2363
rect 8987 2329 8999 2363
rect 9490 2360 9496 2372
rect 8941 2323 8999 2329
rect 9140 2332 9496 2360
rect 5350 2252 5356 2304
rect 5408 2252 5414 2304
rect 6086 2252 6092 2304
rect 6144 2292 6150 2304
rect 6181 2295 6239 2301
rect 6181 2292 6193 2295
rect 6144 2264 6193 2292
rect 6144 2252 6150 2264
rect 6181 2261 6193 2264
rect 6227 2261 6239 2295
rect 6181 2255 6239 2261
rect 8846 2252 8852 2304
rect 8904 2292 8910 2304
rect 9140 2301 9168 2332
rect 9490 2320 9496 2332
rect 9548 2320 9554 2372
rect 9125 2295 9183 2301
rect 9125 2292 9137 2295
rect 8904 2264 9137 2292
rect 8904 2252 8910 2264
rect 9125 2261 9137 2264
rect 9171 2261 9183 2295
rect 9125 2255 9183 2261
rect 9214 2252 9220 2304
rect 9272 2292 9278 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 9272 2264 9321 2292
rect 9272 2252 9278 2264
rect 9309 2261 9321 2264
rect 9355 2292 9367 2295
rect 9398 2292 9404 2304
rect 9355 2264 9404 2292
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 9398 2252 9404 2264
rect 9456 2252 9462 2304
rect 552 2202 11408 2224
rect 552 2150 1755 2202
rect 1807 2150 1819 2202
rect 1871 2150 1883 2202
rect 1935 2150 1947 2202
rect 1999 2150 2011 2202
rect 2063 2150 4469 2202
rect 4521 2150 4533 2202
rect 4585 2150 4597 2202
rect 4649 2150 4661 2202
rect 4713 2150 4725 2202
rect 4777 2150 7183 2202
rect 7235 2150 7247 2202
rect 7299 2150 7311 2202
rect 7363 2150 7375 2202
rect 7427 2150 7439 2202
rect 7491 2150 9897 2202
rect 9949 2150 9961 2202
rect 10013 2150 10025 2202
rect 10077 2150 10089 2202
rect 10141 2150 10153 2202
rect 10205 2150 11408 2202
rect 552 2128 11408 2150
rect 1486 2048 1492 2100
rect 1544 2088 1550 2100
rect 2409 2091 2467 2097
rect 2409 2088 2421 2091
rect 1544 2060 2421 2088
rect 1544 2048 1550 2060
rect 2409 2057 2421 2060
rect 2455 2057 2467 2091
rect 2409 2051 2467 2057
rect 3694 2048 3700 2100
rect 3752 2088 3758 2100
rect 3789 2091 3847 2097
rect 3789 2088 3801 2091
rect 3752 2060 3801 2088
rect 3752 2048 3758 2060
rect 3789 2057 3801 2060
rect 3835 2057 3847 2091
rect 3789 2051 3847 2057
rect 5074 2048 5080 2100
rect 5132 2088 5138 2100
rect 6825 2091 6883 2097
rect 6825 2088 6837 2091
rect 5132 2060 6837 2088
rect 5132 2048 5138 2060
rect 6825 2057 6837 2060
rect 6871 2057 6883 2091
rect 6825 2051 6883 2057
rect 8757 2091 8815 2097
rect 8757 2057 8769 2091
rect 8803 2088 8815 2091
rect 9306 2088 9312 2100
rect 8803 2060 9312 2088
rect 8803 2057 8815 2060
rect 8757 2051 8815 2057
rect 6840 2020 6868 2051
rect 9306 2048 9312 2060
rect 9364 2048 9370 2100
rect 9214 2020 9220 2032
rect 6840 1992 9220 2020
rect 9214 1980 9220 1992
rect 9272 1980 9278 2032
rect 4798 1912 4804 1964
rect 4856 1952 4862 1964
rect 5077 1955 5135 1961
rect 5077 1952 5089 1955
rect 4856 1924 5089 1952
rect 4856 1912 4862 1924
rect 5077 1921 5089 1924
rect 5123 1921 5135 1955
rect 5077 1915 5135 1921
rect 5350 1912 5356 1964
rect 5408 1912 5414 1964
rect 5994 1912 6000 1964
rect 6052 1952 6058 1964
rect 6052 1924 7052 1952
rect 6052 1912 6058 1924
rect 7024 1893 7052 1924
rect 7009 1887 7067 1893
rect 7009 1853 7021 1887
rect 7055 1853 7067 1887
rect 7009 1847 7067 1853
rect 7193 1887 7251 1893
rect 7193 1853 7205 1887
rect 7239 1884 7251 1887
rect 7742 1884 7748 1896
rect 7239 1856 7748 1884
rect 7239 1853 7251 1856
rect 7193 1847 7251 1853
rect 7742 1844 7748 1856
rect 7800 1844 7806 1896
rect 8846 1844 8852 1896
rect 8904 1844 8910 1896
rect 2682 1776 2688 1828
rect 2740 1776 2746 1828
rect 3510 1776 3516 1828
rect 3568 1816 3574 1828
rect 3697 1819 3755 1825
rect 3697 1816 3709 1819
rect 3568 1788 3709 1816
rect 3568 1776 3574 1788
rect 3697 1785 3709 1788
rect 3743 1785 3755 1819
rect 3697 1779 3755 1785
rect 6086 1776 6092 1828
rect 6144 1776 6150 1828
rect 7101 1751 7159 1757
rect 7101 1717 7113 1751
rect 7147 1748 7159 1751
rect 7190 1748 7196 1760
rect 7147 1720 7196 1748
rect 7147 1717 7159 1720
rect 7101 1711 7159 1717
rect 7190 1708 7196 1720
rect 7248 1708 7254 1760
rect 8386 1708 8392 1760
rect 8444 1708 8450 1760
rect 552 1658 11568 1680
rect 552 1606 3112 1658
rect 3164 1606 3176 1658
rect 3228 1606 3240 1658
rect 3292 1606 3304 1658
rect 3356 1606 3368 1658
rect 3420 1606 5826 1658
rect 5878 1606 5890 1658
rect 5942 1606 5954 1658
rect 6006 1606 6018 1658
rect 6070 1606 6082 1658
rect 6134 1606 8540 1658
rect 8592 1606 8604 1658
rect 8656 1606 8668 1658
rect 8720 1606 8732 1658
rect 8784 1606 8796 1658
rect 8848 1606 11254 1658
rect 11306 1606 11318 1658
rect 11370 1606 11382 1658
rect 11434 1606 11446 1658
rect 11498 1606 11510 1658
rect 11562 1606 11568 1658
rect 552 1584 11568 1606
rect 2682 1504 2688 1556
rect 2740 1504 2746 1556
rect 2853 1547 2911 1553
rect 2853 1513 2865 1547
rect 2899 1544 2911 1547
rect 2899 1516 3464 1544
rect 2899 1513 2911 1516
rect 2853 1507 2911 1513
rect 3053 1479 3111 1485
rect 3053 1445 3065 1479
rect 3099 1476 3111 1479
rect 3145 1479 3203 1485
rect 3145 1476 3157 1479
rect 3099 1448 3157 1476
rect 3099 1445 3111 1448
rect 3053 1439 3111 1445
rect 3145 1445 3157 1448
rect 3191 1445 3203 1479
rect 3345 1479 3403 1485
rect 3345 1476 3357 1479
rect 3145 1439 3203 1445
rect 3344 1445 3357 1476
rect 3391 1445 3403 1479
rect 3436 1476 3464 1516
rect 3510 1504 3516 1556
rect 3568 1504 3574 1556
rect 3605 1547 3663 1553
rect 3605 1513 3617 1547
rect 3651 1513 3663 1547
rect 3605 1507 3663 1513
rect 7653 1547 7711 1553
rect 7653 1513 7665 1547
rect 7699 1513 7711 1547
rect 7653 1507 7711 1513
rect 3620 1476 3648 1507
rect 3436 1448 3648 1476
rect 3344 1439 3403 1445
rect 1394 1368 1400 1420
rect 1452 1408 1458 1420
rect 3068 1408 3096 1439
rect 1452 1380 3096 1408
rect 3344 1408 3372 1439
rect 7190 1436 7196 1488
rect 7248 1436 7254 1488
rect 3973 1411 4031 1417
rect 3973 1408 3985 1411
rect 3344 1380 3985 1408
rect 1452 1368 1458 1380
rect 3973 1377 3985 1380
rect 4019 1408 4031 1411
rect 5534 1408 5540 1420
rect 4019 1380 5540 1408
rect 4019 1377 4031 1380
rect 3973 1371 4031 1377
rect 5534 1368 5540 1380
rect 5592 1368 5598 1420
rect 7668 1408 7696 1507
rect 7742 1504 7748 1556
rect 7800 1544 7806 1556
rect 10137 1547 10195 1553
rect 10137 1544 10149 1547
rect 7800 1516 10149 1544
rect 7800 1504 7806 1516
rect 10137 1513 10149 1516
rect 10183 1513 10195 1547
rect 10137 1507 10195 1513
rect 8205 1411 8263 1417
rect 8205 1408 8217 1411
rect 7668 1380 8217 1408
rect 8205 1377 8217 1380
rect 8251 1408 8263 1411
rect 8294 1408 8300 1420
rect 8251 1380 8300 1408
rect 8251 1377 8263 1380
rect 8205 1371 8263 1377
rect 8294 1368 8300 1380
rect 8352 1368 8358 1420
rect 10321 1411 10379 1417
rect 10321 1377 10333 1411
rect 10367 1408 10379 1411
rect 10686 1408 10692 1420
rect 10367 1380 10692 1408
rect 10367 1377 10379 1380
rect 10321 1371 10379 1377
rect 10686 1368 10692 1380
rect 10744 1368 10750 1420
rect 4062 1300 4068 1352
rect 4120 1300 4126 1352
rect 4798 1300 4804 1352
rect 4856 1340 4862 1352
rect 5905 1343 5963 1349
rect 5905 1340 5917 1343
rect 4856 1312 5917 1340
rect 4856 1300 4862 1312
rect 5905 1309 5917 1312
rect 5951 1309 5963 1343
rect 5905 1303 5963 1309
rect 6181 1343 6239 1349
rect 6181 1309 6193 1343
rect 6227 1340 6239 1343
rect 8113 1343 8171 1349
rect 6227 1312 7880 1340
rect 6227 1309 6239 1312
rect 6181 1303 6239 1309
rect 7852 1281 7880 1312
rect 8113 1309 8125 1343
rect 8159 1340 8171 1343
rect 8386 1340 8392 1352
rect 8159 1312 8392 1340
rect 8159 1309 8171 1312
rect 8113 1303 8171 1309
rect 8386 1300 8392 1312
rect 8444 1300 8450 1352
rect 7837 1275 7895 1281
rect 7837 1241 7849 1275
rect 7883 1241 7895 1275
rect 7837 1235 7895 1241
rect 2869 1207 2927 1213
rect 2869 1173 2881 1207
rect 2915 1204 2927 1207
rect 3326 1204 3332 1216
rect 2915 1176 3332 1204
rect 2915 1173 2927 1176
rect 2869 1167 2927 1173
rect 3326 1164 3332 1176
rect 3384 1164 3390 1216
rect 552 1114 11408 1136
rect 552 1062 1755 1114
rect 1807 1062 1819 1114
rect 1871 1062 1883 1114
rect 1935 1062 1947 1114
rect 1999 1062 2011 1114
rect 2063 1062 4469 1114
rect 4521 1062 4533 1114
rect 4585 1062 4597 1114
rect 4649 1062 4661 1114
rect 4713 1062 4725 1114
rect 4777 1062 7183 1114
rect 7235 1062 7247 1114
rect 7299 1062 7311 1114
rect 7363 1062 7375 1114
rect 7427 1062 7439 1114
rect 7491 1062 9897 1114
rect 9949 1062 9961 1114
rect 10013 1062 10025 1114
rect 10077 1062 10089 1114
rect 10141 1062 10153 1114
rect 10205 1062 11408 1114
rect 552 1040 11408 1062
rect 1394 960 1400 1012
rect 1452 960 1458 1012
rect 3326 960 3332 1012
rect 3384 1000 3390 1012
rect 3605 1003 3663 1009
rect 3605 1000 3617 1003
rect 3384 972 3617 1000
rect 3384 960 3390 972
rect 3605 969 3617 972
rect 3651 969 3663 1003
rect 3605 963 3663 969
rect 5534 960 5540 1012
rect 5592 1000 5598 1012
rect 5997 1003 6055 1009
rect 5997 1000 6009 1003
rect 5592 972 6009 1000
rect 5592 960 5598 972
rect 5997 969 6009 972
rect 6043 969 6055 1003
rect 5997 963 6055 969
rect 4062 892 4068 944
rect 4120 932 4126 944
rect 8389 935 8447 941
rect 8389 932 8401 935
rect 4120 904 8401 932
rect 4120 892 4126 904
rect 8389 901 8401 904
rect 8435 901 8447 935
rect 8389 895 8447 901
rect 1118 756 1124 808
rect 1176 796 1182 808
rect 1213 799 1271 805
rect 1213 796 1225 799
rect 1176 768 1225 796
rect 1176 756 1182 768
rect 1213 765 1225 768
rect 1259 765 1271 799
rect 1213 759 1271 765
rect 3510 756 3516 808
rect 3568 796 3574 808
rect 3789 799 3847 805
rect 3789 796 3801 799
rect 3568 768 3801 796
rect 3568 756 3574 768
rect 3789 765 3801 768
rect 3835 765 3847 799
rect 3789 759 3847 765
rect 6178 756 6184 808
rect 6236 756 6242 808
rect 8294 756 8300 808
rect 8352 796 8358 808
rect 8573 799 8631 805
rect 8573 796 8585 799
rect 8352 768 8585 796
rect 8352 756 8358 768
rect 8573 765 8585 768
rect 8619 765 8631 799
rect 8573 759 8631 765
rect 552 570 11568 592
rect 552 518 3112 570
rect 3164 518 3176 570
rect 3228 518 3240 570
rect 3292 518 3304 570
rect 3356 518 3368 570
rect 3420 518 5826 570
rect 5878 518 5890 570
rect 5942 518 5954 570
rect 6006 518 6018 570
rect 6070 518 6082 570
rect 6134 518 8540 570
rect 8592 518 8604 570
rect 8656 518 8668 570
rect 8720 518 8732 570
rect 8784 518 8796 570
rect 8848 518 11254 570
rect 11306 518 11318 570
rect 11370 518 11382 570
rect 11434 518 11446 570
rect 11498 518 11510 570
rect 11562 518 11568 570
rect 552 496 11568 518
<< via1 >>
rect 3112 9222 3164 9274
rect 3176 9222 3228 9274
rect 3240 9222 3292 9274
rect 3304 9222 3356 9274
rect 3368 9222 3420 9274
rect 5826 9222 5878 9274
rect 5890 9222 5942 9274
rect 5954 9222 6006 9274
rect 6018 9222 6070 9274
rect 6082 9222 6134 9274
rect 8540 9222 8592 9274
rect 8604 9222 8656 9274
rect 8668 9222 8720 9274
rect 8732 9222 8784 9274
rect 8796 9222 8848 9274
rect 11254 9222 11306 9274
rect 11318 9222 11370 9274
rect 11382 9222 11434 9274
rect 11446 9222 11498 9274
rect 11510 9222 11562 9274
rect 8300 9120 8352 9172
rect 8668 8916 8720 8968
rect 8944 8891 8996 8900
rect 8944 8857 8953 8891
rect 8953 8857 8987 8891
rect 8987 8857 8996 8891
rect 8944 8848 8996 8857
rect 1755 8678 1807 8730
rect 1819 8678 1871 8730
rect 1883 8678 1935 8730
rect 1947 8678 1999 8730
rect 2011 8678 2063 8730
rect 4469 8678 4521 8730
rect 4533 8678 4585 8730
rect 4597 8678 4649 8730
rect 4661 8678 4713 8730
rect 4725 8678 4777 8730
rect 7183 8678 7235 8730
rect 7247 8678 7299 8730
rect 7311 8678 7363 8730
rect 7375 8678 7427 8730
rect 7439 8678 7491 8730
rect 9897 8678 9949 8730
rect 9961 8678 10013 8730
rect 10025 8678 10077 8730
rect 10089 8678 10141 8730
rect 10153 8678 10205 8730
rect 8576 8576 8628 8628
rect 8944 8576 8996 8628
rect 9404 8576 9456 8628
rect 10692 8619 10744 8628
rect 10692 8585 10701 8619
rect 10701 8585 10735 8619
rect 10735 8585 10744 8619
rect 10692 8576 10744 8585
rect 6736 8508 6788 8560
rect 3424 8372 3476 8424
rect 4804 8372 4856 8424
rect 8668 8440 8720 8492
rect 3608 8347 3660 8356
rect 3608 8313 3642 8347
rect 3642 8313 3660 8347
rect 3608 8304 3660 8313
rect 5632 8347 5684 8356
rect 5632 8313 5666 8347
rect 5666 8313 5684 8347
rect 5632 8304 5684 8313
rect 4712 8279 4764 8288
rect 4712 8245 4721 8279
rect 4721 8245 4755 8279
rect 4755 8245 4764 8279
rect 4712 8236 4764 8245
rect 6184 8236 6236 8288
rect 8116 8415 8168 8424
rect 8116 8381 8125 8415
rect 8125 8381 8159 8415
rect 8159 8381 8168 8415
rect 8116 8372 8168 8381
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 9036 8415 9088 8424
rect 9036 8381 9045 8415
rect 9045 8381 9079 8415
rect 9079 8381 9088 8415
rect 9036 8372 9088 8381
rect 8944 8304 8996 8356
rect 6736 8279 6788 8288
rect 6736 8245 6745 8279
rect 6745 8245 6779 8279
rect 6779 8245 6788 8279
rect 6736 8236 6788 8245
rect 8300 8236 8352 8288
rect 9128 8236 9180 8288
rect 3112 8134 3164 8186
rect 3176 8134 3228 8186
rect 3240 8134 3292 8186
rect 3304 8134 3356 8186
rect 3368 8134 3420 8186
rect 5826 8134 5878 8186
rect 5890 8134 5942 8186
rect 5954 8134 6006 8186
rect 6018 8134 6070 8186
rect 6082 8134 6134 8186
rect 8540 8134 8592 8186
rect 8604 8134 8656 8186
rect 8668 8134 8720 8186
rect 8732 8134 8784 8186
rect 8796 8134 8848 8186
rect 11254 8134 11306 8186
rect 11318 8134 11370 8186
rect 11382 8134 11434 8186
rect 11446 8134 11498 8186
rect 11510 8134 11562 8186
rect 4160 8032 4212 8084
rect 4804 8032 4856 8084
rect 3976 7896 4028 7948
rect 4344 7896 4396 7948
rect 4712 7896 4764 7948
rect 5632 7964 5684 8016
rect 5356 7939 5408 7948
rect 5356 7905 5365 7939
rect 5365 7905 5399 7939
rect 5399 7905 5408 7939
rect 8024 7964 8076 8016
rect 5356 7896 5408 7905
rect 6736 7896 6788 7948
rect 6920 7896 6972 7948
rect 9036 7896 9088 7948
rect 9312 7896 9364 7948
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 3608 7760 3660 7812
rect 4068 7803 4120 7812
rect 4068 7769 4077 7803
rect 4077 7769 4111 7803
rect 4111 7769 4120 7803
rect 4068 7760 4120 7769
rect 6552 7760 6604 7812
rect 7104 7828 7156 7880
rect 8116 7760 8168 7812
rect 7012 7692 7064 7744
rect 8024 7692 8076 7744
rect 8576 7692 8628 7744
rect 9036 7692 9088 7744
rect 10600 7735 10652 7744
rect 10600 7701 10609 7735
rect 10609 7701 10643 7735
rect 10643 7701 10652 7735
rect 10600 7692 10652 7701
rect 1755 7590 1807 7642
rect 1819 7590 1871 7642
rect 1883 7590 1935 7642
rect 1947 7590 1999 7642
rect 2011 7590 2063 7642
rect 4469 7590 4521 7642
rect 4533 7590 4585 7642
rect 4597 7590 4649 7642
rect 4661 7590 4713 7642
rect 4725 7590 4777 7642
rect 7183 7590 7235 7642
rect 7247 7590 7299 7642
rect 7311 7590 7363 7642
rect 7375 7590 7427 7642
rect 7439 7590 7491 7642
rect 9897 7590 9949 7642
rect 9961 7590 10013 7642
rect 10025 7590 10077 7642
rect 10089 7590 10141 7642
rect 10153 7590 10205 7642
rect 4068 7488 4120 7540
rect 4160 7531 4212 7540
rect 4160 7497 4169 7531
rect 4169 7497 4203 7531
rect 4203 7497 4212 7531
rect 4160 7488 4212 7497
rect 6460 7488 6512 7540
rect 6552 7531 6604 7540
rect 6552 7497 6561 7531
rect 6561 7497 6595 7531
rect 6595 7497 6604 7531
rect 6552 7488 6604 7497
rect 8944 7488 8996 7540
rect 9312 7488 9364 7540
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 6368 7352 6420 7404
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 1124 7284 1176 7336
rect 3516 7284 3568 7336
rect 3976 7284 4028 7336
rect 4712 7284 4764 7336
rect 5356 7284 5408 7336
rect 2320 7216 2372 7268
rect 4344 7259 4396 7268
rect 4344 7225 4353 7259
rect 4353 7225 4387 7259
rect 4387 7225 4396 7259
rect 4344 7216 4396 7225
rect 3608 7148 3660 7200
rect 4436 7148 4488 7200
rect 7104 7284 7156 7336
rect 8392 7420 8444 7472
rect 7748 7284 7800 7336
rect 8024 7327 8076 7336
rect 8024 7293 8033 7327
rect 8033 7293 8067 7327
rect 8067 7293 8076 7327
rect 8024 7284 8076 7293
rect 8300 7284 8352 7336
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 9128 7352 9180 7404
rect 10600 7395 10652 7404
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 9404 7284 9456 7336
rect 11060 7327 11112 7336
rect 11060 7293 11069 7327
rect 11069 7293 11103 7327
rect 11103 7293 11112 7327
rect 11060 7284 11112 7293
rect 8116 7148 8168 7200
rect 8208 7148 8260 7200
rect 10876 7191 10928 7200
rect 10876 7157 10885 7191
rect 10885 7157 10919 7191
rect 10919 7157 10928 7191
rect 10876 7148 10928 7157
rect 3112 7046 3164 7098
rect 3176 7046 3228 7098
rect 3240 7046 3292 7098
rect 3304 7046 3356 7098
rect 3368 7046 3420 7098
rect 5826 7046 5878 7098
rect 5890 7046 5942 7098
rect 5954 7046 6006 7098
rect 6018 7046 6070 7098
rect 6082 7046 6134 7098
rect 8540 7046 8592 7098
rect 8604 7046 8656 7098
rect 8668 7046 8720 7098
rect 8732 7046 8784 7098
rect 8796 7046 8848 7098
rect 11254 7046 11306 7098
rect 11318 7046 11370 7098
rect 11382 7046 11434 7098
rect 11446 7046 11498 7098
rect 11510 7046 11562 7098
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 2320 6808 2372 6860
rect 2412 6808 2464 6860
rect 3608 6944 3660 6996
rect 7748 6944 7800 6996
rect 9128 6944 9180 6996
rect 4068 6876 4120 6928
rect 1400 6740 1452 6792
rect 1860 6783 1912 6792
rect 1860 6749 1869 6783
rect 1869 6749 1903 6783
rect 1903 6749 1912 6783
rect 1860 6740 1912 6749
rect 1308 6604 1360 6656
rect 1676 6604 1728 6656
rect 3240 6851 3292 6860
rect 3240 6817 3249 6851
rect 3249 6817 3283 6851
rect 3283 6817 3292 6851
rect 3240 6808 3292 6817
rect 3056 6740 3108 6792
rect 3976 6808 4028 6860
rect 4160 6851 4212 6860
rect 4160 6817 4169 6851
rect 4169 6817 4203 6851
rect 4203 6817 4212 6851
rect 4160 6808 4212 6817
rect 5172 6876 5224 6928
rect 8024 6876 8076 6928
rect 4896 6808 4948 6860
rect 7656 6851 7708 6860
rect 7656 6817 7665 6851
rect 7665 6817 7699 6851
rect 7699 6817 7708 6851
rect 7656 6808 7708 6817
rect 8300 6876 8352 6928
rect 5264 6740 5316 6792
rect 6552 6740 6604 6792
rect 7104 6672 7156 6724
rect 9036 6808 9088 6860
rect 9588 6672 9640 6724
rect 9772 6808 9824 6860
rect 10416 6851 10468 6860
rect 10416 6817 10425 6851
rect 10425 6817 10459 6851
rect 10459 6817 10468 6851
rect 10416 6808 10468 6817
rect 10876 6808 10928 6860
rect 2228 6647 2280 6656
rect 2228 6613 2237 6647
rect 2237 6613 2271 6647
rect 2271 6613 2280 6647
rect 2228 6604 2280 6613
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 4252 6604 4304 6656
rect 8208 6604 8260 6656
rect 8392 6604 8444 6656
rect 9680 6604 9732 6656
rect 1755 6502 1807 6554
rect 1819 6502 1871 6554
rect 1883 6502 1935 6554
rect 1947 6502 1999 6554
rect 2011 6502 2063 6554
rect 4469 6502 4521 6554
rect 4533 6502 4585 6554
rect 4597 6502 4649 6554
rect 4661 6502 4713 6554
rect 4725 6502 4777 6554
rect 7183 6502 7235 6554
rect 7247 6502 7299 6554
rect 7311 6502 7363 6554
rect 7375 6502 7427 6554
rect 7439 6502 7491 6554
rect 9897 6502 9949 6554
rect 9961 6502 10013 6554
rect 10025 6502 10077 6554
rect 10089 6502 10141 6554
rect 10153 6502 10205 6554
rect 1400 6400 1452 6452
rect 2228 6400 2280 6452
rect 3240 6400 3292 6452
rect 3884 6400 3936 6452
rect 4344 6400 4396 6452
rect 5264 6443 5316 6452
rect 5264 6409 5273 6443
rect 5273 6409 5307 6443
rect 5307 6409 5316 6443
rect 5264 6400 5316 6409
rect 5356 6400 5408 6452
rect 6828 6400 6880 6452
rect 7656 6443 7708 6452
rect 7656 6409 7665 6443
rect 7665 6409 7699 6443
rect 7699 6409 7708 6443
rect 7656 6400 7708 6409
rect 2412 6375 2464 6384
rect 2412 6341 2421 6375
rect 2421 6341 2455 6375
rect 2455 6341 2464 6375
rect 2412 6332 2464 6341
rect 2320 6264 2372 6316
rect 3056 6375 3108 6384
rect 3056 6341 3065 6375
rect 3065 6341 3099 6375
rect 3099 6341 3108 6375
rect 3056 6332 3108 6341
rect 4896 6332 4948 6384
rect 1124 6196 1176 6248
rect 1308 6239 1360 6248
rect 1308 6205 1342 6239
rect 1342 6205 1360 6239
rect 1308 6196 1360 6205
rect 5264 6264 5316 6316
rect 5172 6239 5224 6248
rect 5172 6205 5181 6239
rect 5181 6205 5215 6239
rect 5215 6205 5224 6239
rect 5172 6196 5224 6205
rect 3516 6171 3568 6180
rect 3516 6137 3525 6171
rect 3525 6137 3559 6171
rect 3559 6137 3568 6171
rect 3516 6128 3568 6137
rect 6920 6196 6972 6248
rect 8300 6196 8352 6248
rect 7564 6171 7616 6180
rect 7564 6137 7573 6171
rect 7573 6137 7607 6171
rect 7607 6137 7616 6171
rect 7564 6128 7616 6137
rect 8944 6239 8996 6248
rect 8944 6205 8953 6239
rect 8953 6205 8987 6239
rect 8987 6205 8996 6239
rect 8944 6196 8996 6205
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 2872 6060 2924 6112
rect 9680 6128 9732 6180
rect 7840 6060 7892 6112
rect 9772 6060 9824 6112
rect 3112 5958 3164 6010
rect 3176 5958 3228 6010
rect 3240 5958 3292 6010
rect 3304 5958 3356 6010
rect 3368 5958 3420 6010
rect 5826 5958 5878 6010
rect 5890 5958 5942 6010
rect 5954 5958 6006 6010
rect 6018 5958 6070 6010
rect 6082 5958 6134 6010
rect 8540 5958 8592 6010
rect 8604 5958 8656 6010
rect 8668 5958 8720 6010
rect 8732 5958 8784 6010
rect 8796 5958 8848 6010
rect 11254 5958 11306 6010
rect 11318 5958 11370 6010
rect 11382 5958 11434 6010
rect 11446 5958 11498 6010
rect 11510 5958 11562 6010
rect 2136 5856 2188 5908
rect 2596 5856 2648 5908
rect 2964 5856 3016 5908
rect 4896 5899 4948 5908
rect 4896 5865 4905 5899
rect 4905 5865 4939 5899
rect 4939 5865 4948 5899
rect 4896 5856 4948 5865
rect 5172 5856 5224 5908
rect 2412 5788 2464 5840
rect 3976 5788 4028 5840
rect 1676 5720 1728 5772
rect 2780 5720 2832 5772
rect 1308 5652 1360 5704
rect 2872 5652 2924 5704
rect 4804 5720 4856 5772
rect 6552 5899 6604 5908
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 7748 5856 7800 5908
rect 8024 5899 8076 5908
rect 8024 5865 8033 5899
rect 8033 5865 8067 5899
rect 8067 5865 8076 5899
rect 8024 5856 8076 5865
rect 8300 5899 8352 5908
rect 8300 5865 8309 5899
rect 8309 5865 8343 5899
rect 8343 5865 8352 5899
rect 8300 5856 8352 5865
rect 3516 5695 3568 5704
rect 3516 5661 3525 5695
rect 3525 5661 3559 5695
rect 3559 5661 3568 5695
rect 3516 5652 3568 5661
rect 7656 5720 7708 5772
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 7840 5652 7892 5704
rect 8208 5763 8260 5772
rect 8208 5729 8217 5763
rect 8217 5729 8251 5763
rect 8251 5729 8260 5763
rect 8208 5720 8260 5729
rect 9864 5788 9916 5840
rect 9588 5720 9640 5772
rect 3424 5584 3476 5636
rect 1584 5516 1636 5568
rect 3148 5559 3200 5568
rect 3148 5525 3157 5559
rect 3157 5525 3191 5559
rect 3191 5525 3200 5559
rect 3148 5516 3200 5525
rect 4988 5559 5040 5568
rect 4988 5525 4997 5559
rect 4997 5525 5031 5559
rect 5031 5525 5040 5559
rect 4988 5516 5040 5525
rect 8484 5516 8536 5568
rect 9588 5559 9640 5568
rect 9588 5525 9597 5559
rect 9597 5525 9631 5559
rect 9631 5525 9640 5559
rect 9588 5516 9640 5525
rect 1755 5414 1807 5466
rect 1819 5414 1871 5466
rect 1883 5414 1935 5466
rect 1947 5414 1999 5466
rect 2011 5414 2063 5466
rect 4469 5414 4521 5466
rect 4533 5414 4585 5466
rect 4597 5414 4649 5466
rect 4661 5414 4713 5466
rect 4725 5414 4777 5466
rect 7183 5414 7235 5466
rect 7247 5414 7299 5466
rect 7311 5414 7363 5466
rect 7375 5414 7427 5466
rect 7439 5414 7491 5466
rect 9897 5414 9949 5466
rect 9961 5414 10013 5466
rect 10025 5414 10077 5466
rect 10089 5414 10141 5466
rect 10153 5414 10205 5466
rect 2596 5312 2648 5364
rect 4160 5312 4212 5364
rect 4252 5355 4304 5364
rect 4252 5321 4261 5355
rect 4261 5321 4295 5355
rect 4295 5321 4304 5355
rect 4252 5312 4304 5321
rect 2872 5244 2924 5296
rect 2228 5176 2280 5228
rect 9496 5312 9548 5364
rect 6368 5244 6420 5296
rect 2780 5108 2832 5160
rect 3148 5108 3200 5160
rect 3424 5108 3476 5160
rect 3608 5108 3660 5160
rect 7656 5176 7708 5228
rect 7748 5151 7800 5160
rect 7748 5117 7752 5151
rect 7752 5117 7786 5151
rect 7786 5117 7800 5151
rect 3884 5040 3936 5092
rect 4712 5040 4764 5092
rect 6184 5040 6236 5092
rect 6920 5040 6972 5092
rect 7748 5108 7800 5117
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 8300 5108 8352 5160
rect 8392 5108 8444 5160
rect 10416 5108 10468 5160
rect 8116 5083 8168 5092
rect 8116 5049 8125 5083
rect 8125 5049 8159 5083
rect 8159 5049 8168 5083
rect 8116 5040 8168 5049
rect 9588 5040 9640 5092
rect 1400 4972 1452 5024
rect 2780 4972 2832 5024
rect 4988 4972 5040 5024
rect 6828 4972 6880 5024
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 7472 5015 7524 5024
rect 7472 4981 7481 5015
rect 7481 4981 7515 5015
rect 7515 4981 7524 5015
rect 7472 4972 7524 4981
rect 10232 4972 10284 5024
rect 3112 4870 3164 4922
rect 3176 4870 3228 4922
rect 3240 4870 3292 4922
rect 3304 4870 3356 4922
rect 3368 4870 3420 4922
rect 5826 4870 5878 4922
rect 5890 4870 5942 4922
rect 5954 4870 6006 4922
rect 6018 4870 6070 4922
rect 6082 4870 6134 4922
rect 8540 4870 8592 4922
rect 8604 4870 8656 4922
rect 8668 4870 8720 4922
rect 8732 4870 8784 4922
rect 8796 4870 8848 4922
rect 11254 4870 11306 4922
rect 11318 4870 11370 4922
rect 11382 4870 11434 4922
rect 11446 4870 11498 4922
rect 11510 4870 11562 4922
rect 1308 4768 1360 4820
rect 2228 4768 2280 4820
rect 2780 4811 2832 4820
rect 2780 4777 2789 4811
rect 2789 4777 2823 4811
rect 2823 4777 2832 4811
rect 2780 4768 2832 4777
rect 6184 4768 6236 4820
rect 7472 4768 7524 4820
rect 8116 4768 8168 4820
rect 1400 4700 1452 4752
rect 1584 4743 1636 4752
rect 1584 4709 1618 4743
rect 1618 4709 1636 4743
rect 1584 4700 1636 4709
rect 2596 4700 2648 4752
rect 3792 4700 3844 4752
rect 1124 4564 1176 4616
rect 3884 4675 3936 4684
rect 3884 4641 3893 4675
rect 3893 4641 3927 4675
rect 3927 4641 3936 4675
rect 3884 4632 3936 4641
rect 7012 4700 7064 4752
rect 10232 4700 10284 4752
rect 6368 4632 6420 4684
rect 6828 4675 6880 4684
rect 6828 4641 6837 4675
rect 6837 4641 6871 4675
rect 6871 4641 6880 4675
rect 6828 4632 6880 4641
rect 9128 4632 9180 4684
rect 1676 4428 1728 4480
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 9680 4564 9732 4616
rect 1755 4326 1807 4378
rect 1819 4326 1871 4378
rect 1883 4326 1935 4378
rect 1947 4326 1999 4378
rect 2011 4326 2063 4378
rect 4469 4326 4521 4378
rect 4533 4326 4585 4378
rect 4597 4326 4649 4378
rect 4661 4326 4713 4378
rect 4725 4326 4777 4378
rect 7183 4326 7235 4378
rect 7247 4326 7299 4378
rect 7311 4326 7363 4378
rect 7375 4326 7427 4378
rect 7439 4326 7491 4378
rect 9897 4326 9949 4378
rect 9961 4326 10013 4378
rect 10025 4326 10077 4378
rect 10089 4326 10141 4378
rect 10153 4326 10205 4378
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 7748 4224 7800 4276
rect 9772 4267 9824 4276
rect 9772 4233 9781 4267
rect 9781 4233 9815 4267
rect 9815 4233 9824 4267
rect 9772 4224 9824 4233
rect 7656 4199 7708 4208
rect 7656 4165 7665 4199
rect 7665 4165 7699 4199
rect 7699 4165 7708 4199
rect 7656 4156 7708 4165
rect 3976 4088 4028 4140
rect 2964 4020 3016 4072
rect 3516 4020 3568 4072
rect 4252 4020 4304 4072
rect 5632 4020 5684 4072
rect 6368 4020 6420 4072
rect 8300 4088 8352 4140
rect 8944 4088 8996 4140
rect 9588 4131 9640 4140
rect 9588 4097 9597 4131
rect 9597 4097 9631 4131
rect 9631 4097 9640 4131
rect 9588 4088 9640 4097
rect 7748 4020 7800 4072
rect 2872 3952 2924 4004
rect 7932 4020 7984 4072
rect 8116 4063 8168 4072
rect 8116 4029 8125 4063
rect 8125 4029 8159 4063
rect 8159 4029 8168 4063
rect 8116 4020 8168 4029
rect 8208 4020 8260 4072
rect 8760 4020 8812 4072
rect 9036 4063 9088 4072
rect 9036 4029 9045 4063
rect 9045 4029 9079 4063
rect 9079 4029 9088 4063
rect 9036 4020 9088 4029
rect 9128 4063 9180 4072
rect 9128 4029 9137 4063
rect 9137 4029 9171 4063
rect 9171 4029 9180 4063
rect 9128 4020 9180 4029
rect 9312 4020 9364 4072
rect 9772 4020 9824 4072
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 6184 3884 6236 3936
rect 6920 3884 6972 3936
rect 8024 3927 8076 3936
rect 8024 3893 8033 3927
rect 8033 3893 8067 3927
rect 8067 3893 8076 3927
rect 8024 3884 8076 3893
rect 3112 3782 3164 3834
rect 3176 3782 3228 3834
rect 3240 3782 3292 3834
rect 3304 3782 3356 3834
rect 3368 3782 3420 3834
rect 5826 3782 5878 3834
rect 5890 3782 5942 3834
rect 5954 3782 6006 3834
rect 6018 3782 6070 3834
rect 6082 3782 6134 3834
rect 8540 3782 8592 3834
rect 8604 3782 8656 3834
rect 8668 3782 8720 3834
rect 8732 3782 8784 3834
rect 8796 3782 8848 3834
rect 11254 3782 11306 3834
rect 11318 3782 11370 3834
rect 11382 3782 11434 3834
rect 11446 3782 11498 3834
rect 11510 3782 11562 3834
rect 3792 3680 3844 3732
rect 8116 3680 8168 3732
rect 9036 3680 9088 3732
rect 2964 3612 3016 3664
rect 2596 3587 2648 3596
rect 2596 3553 2630 3587
rect 2630 3553 2648 3587
rect 2596 3544 2648 3553
rect 5724 3544 5776 3596
rect 6644 3587 6696 3596
rect 6644 3553 6653 3587
rect 6653 3553 6687 3587
rect 6687 3553 6696 3587
rect 6644 3544 6696 3553
rect 4896 3340 4948 3392
rect 7748 3587 7800 3596
rect 7748 3553 7757 3587
rect 7757 3553 7791 3587
rect 7791 3553 7800 3587
rect 7748 3544 7800 3553
rect 7932 3587 7984 3596
rect 7932 3553 7941 3587
rect 7941 3553 7975 3587
rect 7975 3553 7984 3587
rect 7932 3544 7984 3553
rect 8392 3655 8444 3664
rect 8392 3621 8401 3655
rect 8401 3621 8435 3655
rect 8435 3621 8444 3655
rect 8392 3612 8444 3621
rect 8208 3544 8260 3596
rect 8484 3544 8536 3596
rect 9036 3544 9088 3596
rect 9312 3587 9364 3596
rect 9312 3553 9321 3587
rect 9321 3553 9355 3587
rect 9355 3553 9364 3587
rect 9312 3544 9364 3553
rect 8300 3476 8352 3528
rect 8576 3476 8628 3528
rect 9128 3476 9180 3528
rect 9588 3587 9640 3596
rect 9588 3553 9597 3587
rect 9597 3553 9631 3587
rect 9631 3553 9640 3587
rect 9588 3544 9640 3553
rect 10232 3587 10284 3596
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 10416 3476 10468 3528
rect 7932 3340 7984 3392
rect 9404 3340 9456 3392
rect 1755 3238 1807 3290
rect 1819 3238 1871 3290
rect 1883 3238 1935 3290
rect 1947 3238 1999 3290
rect 2011 3238 2063 3290
rect 4469 3238 4521 3290
rect 4533 3238 4585 3290
rect 4597 3238 4649 3290
rect 4661 3238 4713 3290
rect 4725 3238 4777 3290
rect 7183 3238 7235 3290
rect 7247 3238 7299 3290
rect 7311 3238 7363 3290
rect 7375 3238 7427 3290
rect 7439 3238 7491 3290
rect 9897 3238 9949 3290
rect 9961 3238 10013 3290
rect 10025 3238 10077 3290
rect 10089 3238 10141 3290
rect 10153 3238 10205 3290
rect 2596 3136 2648 3188
rect 3608 3136 3660 3188
rect 7748 3136 7800 3188
rect 8484 3136 8536 3188
rect 9404 3136 9456 3188
rect 8208 3068 8260 3120
rect 8852 3068 8904 3120
rect 9496 3068 9548 3120
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 9864 3179 9916 3188
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 9864 3136 9916 3145
rect 10416 3179 10468 3188
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 3792 3000 3844 3009
rect 4896 3043 4948 3052
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 3976 2864 4028 2916
rect 6184 2932 6236 2984
rect 8484 3000 8536 3052
rect 9128 3000 9180 3052
rect 6644 2932 6696 2984
rect 8392 2932 8444 2984
rect 4804 2864 4856 2916
rect 8300 2864 8352 2916
rect 8852 2975 8904 2984
rect 8852 2941 8861 2975
rect 8861 2941 8895 2975
rect 8895 2941 8904 2975
rect 8852 2932 8904 2941
rect 9036 2932 9088 2984
rect 9680 2864 9732 2916
rect 8760 2796 8812 2848
rect 9128 2796 9180 2848
rect 9404 2839 9456 2848
rect 9404 2805 9413 2839
rect 9413 2805 9447 2839
rect 9447 2805 9456 2839
rect 9404 2796 9456 2805
rect 9496 2796 9548 2848
rect 3112 2694 3164 2746
rect 3176 2694 3228 2746
rect 3240 2694 3292 2746
rect 3304 2694 3356 2746
rect 3368 2694 3420 2746
rect 5826 2694 5878 2746
rect 5890 2694 5942 2746
rect 5954 2694 6006 2746
rect 6018 2694 6070 2746
rect 6082 2694 6134 2746
rect 8540 2694 8592 2746
rect 8604 2694 8656 2746
rect 8668 2694 8720 2746
rect 8732 2694 8784 2746
rect 8796 2694 8848 2746
rect 11254 2694 11306 2746
rect 11318 2694 11370 2746
rect 11382 2694 11434 2746
rect 11446 2694 11498 2746
rect 11510 2694 11562 2746
rect 6368 2592 6420 2644
rect 7748 2592 7800 2644
rect 9036 2635 9088 2644
rect 9036 2601 9045 2635
rect 9045 2601 9079 2635
rect 9079 2601 9088 2635
rect 9036 2592 9088 2601
rect 5080 2499 5132 2508
rect 5080 2465 5089 2499
rect 5089 2465 5123 2499
rect 5123 2465 5132 2499
rect 5080 2456 5132 2465
rect 5632 2456 5684 2508
rect 6000 2499 6052 2508
rect 6000 2465 6009 2499
rect 6009 2465 6043 2499
rect 6043 2465 6052 2499
rect 6000 2456 6052 2465
rect 8300 2524 8352 2576
rect 8392 2524 8444 2576
rect 9864 2592 9916 2644
rect 5724 2388 5776 2440
rect 8300 2388 8352 2440
rect 9128 2456 9180 2508
rect 5356 2295 5408 2304
rect 5356 2261 5365 2295
rect 5365 2261 5399 2295
rect 5399 2261 5408 2295
rect 5356 2252 5408 2261
rect 6092 2252 6144 2304
rect 8852 2252 8904 2304
rect 9496 2320 9548 2372
rect 9220 2252 9272 2304
rect 9404 2252 9456 2304
rect 1755 2150 1807 2202
rect 1819 2150 1871 2202
rect 1883 2150 1935 2202
rect 1947 2150 1999 2202
rect 2011 2150 2063 2202
rect 4469 2150 4521 2202
rect 4533 2150 4585 2202
rect 4597 2150 4649 2202
rect 4661 2150 4713 2202
rect 4725 2150 4777 2202
rect 7183 2150 7235 2202
rect 7247 2150 7299 2202
rect 7311 2150 7363 2202
rect 7375 2150 7427 2202
rect 7439 2150 7491 2202
rect 9897 2150 9949 2202
rect 9961 2150 10013 2202
rect 10025 2150 10077 2202
rect 10089 2150 10141 2202
rect 10153 2150 10205 2202
rect 1492 2048 1544 2100
rect 3700 2048 3752 2100
rect 5080 2048 5132 2100
rect 9312 2048 9364 2100
rect 9220 1980 9272 2032
rect 4804 1912 4856 1964
rect 5356 1955 5408 1964
rect 5356 1921 5365 1955
rect 5365 1921 5399 1955
rect 5399 1921 5408 1955
rect 5356 1912 5408 1921
rect 6000 1912 6052 1964
rect 7748 1844 7800 1896
rect 8852 1887 8904 1896
rect 8852 1853 8861 1887
rect 8861 1853 8895 1887
rect 8895 1853 8904 1887
rect 8852 1844 8904 1853
rect 2688 1819 2740 1828
rect 2688 1785 2697 1819
rect 2697 1785 2731 1819
rect 2731 1785 2740 1819
rect 2688 1776 2740 1785
rect 3516 1776 3568 1828
rect 6092 1776 6144 1828
rect 7196 1708 7248 1760
rect 8392 1751 8444 1760
rect 8392 1717 8401 1751
rect 8401 1717 8435 1751
rect 8435 1717 8444 1751
rect 8392 1708 8444 1717
rect 3112 1606 3164 1658
rect 3176 1606 3228 1658
rect 3240 1606 3292 1658
rect 3304 1606 3356 1658
rect 3368 1606 3420 1658
rect 5826 1606 5878 1658
rect 5890 1606 5942 1658
rect 5954 1606 6006 1658
rect 6018 1606 6070 1658
rect 6082 1606 6134 1658
rect 8540 1606 8592 1658
rect 8604 1606 8656 1658
rect 8668 1606 8720 1658
rect 8732 1606 8784 1658
rect 8796 1606 8848 1658
rect 11254 1606 11306 1658
rect 11318 1606 11370 1658
rect 11382 1606 11434 1658
rect 11446 1606 11498 1658
rect 11510 1606 11562 1658
rect 2688 1547 2740 1556
rect 2688 1513 2697 1547
rect 2697 1513 2731 1547
rect 2731 1513 2740 1547
rect 2688 1504 2740 1513
rect 3516 1547 3568 1556
rect 3516 1513 3525 1547
rect 3525 1513 3559 1547
rect 3559 1513 3568 1547
rect 3516 1504 3568 1513
rect 1400 1368 1452 1420
rect 7196 1436 7248 1488
rect 5540 1368 5592 1420
rect 7748 1504 7800 1556
rect 8300 1368 8352 1420
rect 10692 1368 10744 1420
rect 4068 1343 4120 1352
rect 4068 1309 4077 1343
rect 4077 1309 4111 1343
rect 4111 1309 4120 1343
rect 4068 1300 4120 1309
rect 4804 1300 4856 1352
rect 8392 1300 8444 1352
rect 3332 1207 3384 1216
rect 3332 1173 3341 1207
rect 3341 1173 3375 1207
rect 3375 1173 3384 1207
rect 3332 1164 3384 1173
rect 1755 1062 1807 1114
rect 1819 1062 1871 1114
rect 1883 1062 1935 1114
rect 1947 1062 1999 1114
rect 2011 1062 2063 1114
rect 4469 1062 4521 1114
rect 4533 1062 4585 1114
rect 4597 1062 4649 1114
rect 4661 1062 4713 1114
rect 4725 1062 4777 1114
rect 7183 1062 7235 1114
rect 7247 1062 7299 1114
rect 7311 1062 7363 1114
rect 7375 1062 7427 1114
rect 7439 1062 7491 1114
rect 9897 1062 9949 1114
rect 9961 1062 10013 1114
rect 10025 1062 10077 1114
rect 10089 1062 10141 1114
rect 10153 1062 10205 1114
rect 1400 1003 1452 1012
rect 1400 969 1409 1003
rect 1409 969 1443 1003
rect 1443 969 1452 1003
rect 1400 960 1452 969
rect 3332 960 3384 1012
rect 5540 960 5592 1012
rect 4068 892 4120 944
rect 1124 756 1176 808
rect 3516 756 3568 808
rect 6184 799 6236 808
rect 6184 765 6193 799
rect 6193 765 6227 799
rect 6227 765 6236 799
rect 6184 756 6236 765
rect 8300 756 8352 808
rect 3112 518 3164 570
rect 3176 518 3228 570
rect 3240 518 3292 570
rect 3304 518 3356 570
rect 3368 518 3420 570
rect 5826 518 5878 570
rect 5890 518 5942 570
rect 5954 518 6006 570
rect 6018 518 6070 570
rect 6082 518 6134 570
rect 8540 518 8592 570
rect 8604 518 8656 570
rect 8668 518 8720 570
rect 8732 518 8784 570
rect 8796 518 8848 570
rect 11254 518 11306 570
rect 11318 518 11370 570
rect 11382 518 11434 570
rect 11446 518 11498 570
rect 11510 518 11562 570
<< metal2 >>
rect 1122 9738 1178 10000
rect 3514 9738 3570 10000
rect 5906 9738 5962 10000
rect 1122 9710 1348 9738
rect 1122 9600 1178 9710
rect 1124 7336 1176 7342
rect 1124 7278 1176 7284
rect 1136 6254 1164 7278
rect 1320 6914 1348 9710
rect 3514 9710 3740 9738
rect 3514 9600 3570 9710
rect 3112 9276 3420 9285
rect 3112 9274 3118 9276
rect 3174 9274 3198 9276
rect 3254 9274 3278 9276
rect 3334 9274 3358 9276
rect 3414 9274 3420 9276
rect 3174 9222 3176 9274
rect 3356 9222 3358 9274
rect 3112 9220 3118 9222
rect 3174 9220 3198 9222
rect 3254 9220 3278 9222
rect 3334 9220 3358 9222
rect 3414 9220 3420 9222
rect 3112 9211 3420 9220
rect 1755 8732 2063 8741
rect 1755 8730 1761 8732
rect 1817 8730 1841 8732
rect 1897 8730 1921 8732
rect 1977 8730 2001 8732
rect 2057 8730 2063 8732
rect 1817 8678 1819 8730
rect 1999 8678 2001 8730
rect 1755 8676 1761 8678
rect 1817 8676 1841 8678
rect 1897 8676 1921 8678
rect 1977 8676 2001 8678
rect 2057 8676 2063 8678
rect 1755 8667 2063 8676
rect 3424 8424 3476 8430
rect 3476 8372 3556 8378
rect 3424 8366 3556 8372
rect 3436 8350 3556 8366
rect 3112 8188 3420 8197
rect 3112 8186 3118 8188
rect 3174 8186 3198 8188
rect 3254 8186 3278 8188
rect 3334 8186 3358 8188
rect 3414 8186 3420 8188
rect 3174 8134 3176 8186
rect 3356 8134 3358 8186
rect 3112 8132 3118 8134
rect 3174 8132 3198 8134
rect 3254 8132 3278 8134
rect 3334 8132 3358 8134
rect 3414 8132 3420 8134
rect 3112 8123 3420 8132
rect 1755 7644 2063 7653
rect 1755 7642 1761 7644
rect 1817 7642 1841 7644
rect 1897 7642 1921 7644
rect 1977 7642 2001 7644
rect 2057 7642 2063 7644
rect 1817 7590 1819 7642
rect 1999 7590 2001 7642
rect 1755 7588 1761 7590
rect 1817 7588 1841 7590
rect 1897 7588 1921 7590
rect 1977 7588 2001 7590
rect 2057 7588 2063 7590
rect 1755 7579 2063 7588
rect 3528 7342 3556 8350
rect 3608 8356 3660 8362
rect 3608 8298 3660 8304
rect 3620 7818 3648 8298
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2332 7002 2360 7210
rect 3112 7100 3420 7109
rect 3112 7098 3118 7100
rect 3174 7098 3198 7100
rect 3254 7098 3278 7100
rect 3334 7098 3358 7100
rect 3414 7098 3420 7100
rect 3174 7046 3176 7098
rect 3356 7046 3358 7098
rect 3112 7044 3118 7046
rect 3174 7044 3198 7046
rect 3254 7044 3278 7046
rect 3334 7044 3358 7046
rect 3414 7044 3420 7046
rect 3112 7035 3420 7044
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 1320 6886 1532 6914
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1308 6656 1360 6662
rect 1308 6598 1360 6604
rect 1320 6254 1348 6598
rect 1412 6458 1440 6734
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1124 6248 1176 6254
rect 1124 6190 1176 6196
rect 1308 6248 1360 6254
rect 1308 6190 1360 6196
rect 1136 4622 1164 6190
rect 1308 5704 1360 5710
rect 1308 5646 1360 5652
rect 1320 4826 1348 5646
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1308 4820 1360 4826
rect 1308 4762 1360 4768
rect 1412 4758 1440 4966
rect 1400 4752 1452 4758
rect 1400 4694 1452 4700
rect 1124 4616 1176 4622
rect 1124 4558 1176 4564
rect 1504 2106 1532 6886
rect 2424 6866 2636 6882
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2412 6860 2636 6866
rect 2464 6854 2636 6860
rect 2412 6802 2464 6808
rect 1860 6792 1912 6798
rect 1912 6740 2176 6746
rect 1860 6734 2176 6740
rect 1872 6718 2176 6734
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1688 5778 1716 6598
rect 1755 6556 2063 6565
rect 1755 6554 1761 6556
rect 1817 6554 1841 6556
rect 1897 6554 1921 6556
rect 1977 6554 2001 6556
rect 2057 6554 2063 6556
rect 1817 6502 1819 6554
rect 1999 6502 2001 6554
rect 1755 6500 1761 6502
rect 1817 6500 1841 6502
rect 1897 6500 1921 6502
rect 1977 6500 2001 6502
rect 2057 6500 2063 6502
rect 1755 6491 2063 6500
rect 2148 5914 2176 6718
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2240 6458 2268 6598
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2332 6322 2360 6802
rect 2412 6384 2464 6390
rect 2412 6326 2464 6332
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1596 4758 1624 5510
rect 1584 4752 1636 4758
rect 1584 4694 1636 4700
rect 1688 4486 1716 5714
rect 1755 5468 2063 5477
rect 1755 5466 1761 5468
rect 1817 5466 1841 5468
rect 1897 5466 1921 5468
rect 1977 5466 2001 5468
rect 2057 5466 2063 5468
rect 1817 5414 1819 5466
rect 1999 5414 2001 5466
rect 1755 5412 1761 5414
rect 1817 5412 1841 5414
rect 1897 5412 1921 5414
rect 1977 5412 2001 5414
rect 2057 5412 2063 5414
rect 1755 5403 2063 5412
rect 2148 5250 2176 5850
rect 2424 5846 2452 6326
rect 2608 5914 2636 6854
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 3068 6390 3096 6734
rect 3252 6458 3280 6802
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 3068 6202 3096 6326
rect 2976 6174 3096 6202
rect 3528 6186 3556 7278
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3620 7002 3648 7142
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3516 6180 3568 6186
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 2608 5370 2636 5850
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2148 5234 2268 5250
rect 2148 5228 2280 5234
rect 2148 5222 2228 5228
rect 2228 5170 2280 5176
rect 2240 4826 2268 5170
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2608 4758 2636 5306
rect 2792 5166 2820 5714
rect 2884 5710 2912 6054
rect 2976 5914 3004 6174
rect 3516 6122 3568 6128
rect 3112 6012 3420 6021
rect 3112 6010 3118 6012
rect 3174 6010 3198 6012
rect 3254 6010 3278 6012
rect 3334 6010 3358 6012
rect 3414 6010 3420 6012
rect 3174 5958 3176 6010
rect 3356 5958 3358 6010
rect 3112 5956 3118 5958
rect 3174 5956 3198 5958
rect 3254 5956 3278 5958
rect 3334 5956 3358 5958
rect 3414 5956 3420 5958
rect 3112 5947 3420 5956
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 3528 5710 3556 6122
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2792 5030 2820 5102
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 4826 2820 4966
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2596 4752 2648 4758
rect 2596 4694 2648 4700
rect 1676 4480 1728 4486
rect 1676 4422 1728 4428
rect 1688 4282 1716 4422
rect 1755 4380 2063 4389
rect 1755 4378 1761 4380
rect 1817 4378 1841 4380
rect 1897 4378 1921 4380
rect 1977 4378 2001 4380
rect 2057 4378 2063 4380
rect 1817 4326 1819 4378
rect 1999 4326 2001 4378
rect 1755 4324 1761 4326
rect 1817 4324 1841 4326
rect 1897 4324 1921 4326
rect 1977 4324 2001 4326
rect 2057 4324 2063 4326
rect 1755 4315 2063 4324
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 2884 4010 2912 5238
rect 3160 5166 3188 5510
rect 3436 5166 3464 5578
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3112 4924 3420 4933
rect 3112 4922 3118 4924
rect 3174 4922 3198 4924
rect 3254 4922 3278 4924
rect 3334 4922 3358 4924
rect 3414 4922 3420 4924
rect 3174 4870 3176 4922
rect 3356 4870 3358 4922
rect 3112 4868 3118 4870
rect 3174 4868 3198 4870
rect 3254 4868 3278 4870
rect 3334 4868 3358 4870
rect 3414 4868 3420 4870
rect 3112 4859 3420 4868
rect 3528 4078 3556 5646
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2976 3670 3004 4014
rect 3112 3836 3420 3845
rect 3112 3834 3118 3836
rect 3174 3834 3198 3836
rect 3254 3834 3278 3836
rect 3334 3834 3358 3836
rect 3414 3834 3420 3836
rect 3174 3782 3176 3834
rect 3356 3782 3358 3834
rect 3112 3780 3118 3782
rect 3174 3780 3198 3782
rect 3254 3780 3278 3782
rect 3334 3780 3358 3782
rect 3414 3780 3420 3782
rect 3112 3771 3420 3780
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 2596 3596 2648 3602
rect 2596 3538 2648 3544
rect 1755 3292 2063 3301
rect 1755 3290 1761 3292
rect 1817 3290 1841 3292
rect 1897 3290 1921 3292
rect 1977 3290 2001 3292
rect 2057 3290 2063 3292
rect 1817 3238 1819 3290
rect 1999 3238 2001 3290
rect 1755 3236 1761 3238
rect 1817 3236 1841 3238
rect 1897 3236 1921 3238
rect 1977 3236 2001 3238
rect 2057 3236 2063 3238
rect 1755 3227 2063 3236
rect 2608 3194 2636 3538
rect 3620 3194 3648 5102
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3112 2748 3420 2757
rect 3112 2746 3118 2748
rect 3174 2746 3198 2748
rect 3254 2746 3278 2748
rect 3334 2746 3358 2748
rect 3414 2746 3420 2748
rect 3174 2694 3176 2746
rect 3356 2694 3358 2746
rect 3112 2692 3118 2694
rect 3174 2692 3198 2694
rect 3254 2692 3278 2694
rect 3334 2692 3358 2694
rect 3414 2692 3420 2694
rect 3112 2683 3420 2692
rect 1755 2204 2063 2213
rect 1755 2202 1761 2204
rect 1817 2202 1841 2204
rect 1897 2202 1921 2204
rect 1977 2202 2001 2204
rect 2057 2202 2063 2204
rect 1817 2150 1819 2202
rect 1999 2150 2001 2202
rect 1755 2148 1761 2150
rect 1817 2148 1841 2150
rect 1897 2148 1921 2150
rect 1977 2148 2001 2150
rect 2057 2148 2063 2150
rect 1755 2139 2063 2148
rect 3712 2106 3740 9710
rect 5906 9710 6224 9738
rect 5906 9600 5962 9710
rect 5826 9276 6134 9285
rect 5826 9274 5832 9276
rect 5888 9274 5912 9276
rect 5968 9274 5992 9276
rect 6048 9274 6072 9276
rect 6128 9274 6134 9276
rect 5888 9222 5890 9274
rect 6070 9222 6072 9274
rect 5826 9220 5832 9222
rect 5888 9220 5912 9222
rect 5968 9220 5992 9222
rect 6048 9220 6072 9222
rect 6128 9220 6134 9222
rect 5826 9211 6134 9220
rect 4469 8732 4777 8741
rect 4469 8730 4475 8732
rect 4531 8730 4555 8732
rect 4611 8730 4635 8732
rect 4691 8730 4715 8732
rect 4771 8730 4777 8732
rect 4531 8678 4533 8730
rect 4713 8678 4715 8730
rect 4469 8676 4475 8678
rect 4531 8676 4555 8678
rect 4611 8676 4635 8678
rect 4691 8676 4715 8678
rect 4771 8676 4777 8678
rect 4469 8667 4777 8676
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 3988 7342 4016 7890
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 4080 7546 4108 7754
rect 4172 7546 4200 8026
rect 4724 7954 4752 8230
rect 4816 8090 4844 8366
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3976 7336 4028 7342
rect 3976 7278 4028 7284
rect 3988 6866 4016 7278
rect 4080 6934 4108 7482
rect 4356 7274 4384 7890
rect 4469 7644 4777 7653
rect 4469 7642 4475 7644
rect 4531 7642 4555 7644
rect 4611 7642 4635 7644
rect 4691 7642 4715 7644
rect 4771 7642 4777 7644
rect 4531 7590 4533 7642
rect 4713 7590 4715 7642
rect 4469 7588 4475 7590
rect 4531 7588 4555 7590
rect 4611 7588 4635 7590
rect 4691 7588 4715 7590
rect 4771 7588 4777 7590
rect 4469 7579 4777 7588
rect 4816 7410 4844 8026
rect 5644 8022 5672 8298
rect 6196 8294 6224 9710
rect 8298 9600 8354 10000
rect 10690 9600 10746 10000
rect 8312 9178 8340 9600
rect 8540 9276 8848 9285
rect 8540 9274 8546 9276
rect 8602 9274 8626 9276
rect 8682 9274 8706 9276
rect 8762 9274 8786 9276
rect 8842 9274 8848 9276
rect 8602 9222 8604 9274
rect 8784 9222 8786 9274
rect 8540 9220 8546 9222
rect 8602 9220 8626 9222
rect 8682 9220 8706 9222
rect 8762 9220 8786 9222
rect 8842 9220 8848 9222
rect 8540 9211 8848 9220
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 7183 8732 7491 8741
rect 7183 8730 7189 8732
rect 7245 8730 7269 8732
rect 7325 8730 7349 8732
rect 7405 8730 7429 8732
rect 7485 8730 7491 8732
rect 7245 8678 7247 8730
rect 7427 8678 7429 8730
rect 7183 8676 7189 8678
rect 7245 8676 7269 8678
rect 7325 8676 7349 8678
rect 7405 8676 7429 8678
rect 7485 8676 7491 8678
rect 7183 8667 7491 8676
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6748 8294 6776 8502
rect 8588 8430 8616 8570
rect 8680 8498 8708 8910
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8956 8634 8984 8842
rect 9897 8732 10205 8741
rect 9897 8730 9903 8732
rect 9959 8730 9983 8732
rect 10039 8730 10063 8732
rect 10119 8730 10143 8732
rect 10199 8730 10205 8732
rect 9959 8678 9961 8730
rect 10141 8678 10143 8730
rect 9897 8676 9903 8678
rect 9959 8676 9983 8678
rect 10039 8676 10063 8678
rect 10119 8676 10143 8678
rect 10199 8676 10205 8678
rect 9897 8667 10205 8676
rect 10704 8634 10732 9600
rect 11254 9276 11562 9285
rect 11254 9274 11260 9276
rect 11316 9274 11340 9276
rect 11396 9274 11420 9276
rect 11476 9274 11500 9276
rect 11556 9274 11562 9276
rect 11316 9222 11318 9274
rect 11498 9222 11500 9274
rect 11254 9220 11260 9222
rect 11316 9220 11340 9222
rect 11396 9220 11420 9222
rect 11476 9220 11500 9222
rect 11556 9220 11562 9222
rect 11254 9211 11562 9220
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 5826 8188 6134 8197
rect 5826 8186 5832 8188
rect 5888 8186 5912 8188
rect 5968 8186 5992 8188
rect 6048 8186 6072 8188
rect 6128 8186 6134 8188
rect 5888 8134 5890 8186
rect 6070 8134 6072 8186
rect 5826 8132 5832 8134
rect 5888 8132 5912 8134
rect 5968 8132 5992 8134
rect 6048 8132 6072 8134
rect 6128 8132 6134 8134
rect 5826 8123 6134 8132
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 6748 7954 6776 8230
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 5368 7342 5396 7890
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6380 7410 6408 7822
rect 6472 7546 6500 7822
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6564 7546 6592 7754
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 4344 7268 4396 7274
rect 4344 7210 4396 7216
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4068 6928 4120 6934
rect 4448 6914 4476 7142
rect 4068 6870 4120 6876
rect 4356 6886 4476 6914
rect 4724 6914 4752 7278
rect 5826 7100 6134 7109
rect 5826 7098 5832 7100
rect 5888 7098 5912 7100
rect 5968 7098 5992 7100
rect 6048 7098 6072 7100
rect 6128 7098 6134 7100
rect 5888 7046 5890 7098
rect 6070 7046 6072 7098
rect 5826 7044 5832 7046
rect 5888 7044 5912 7046
rect 5968 7044 5992 7046
rect 6048 7044 6072 7046
rect 6128 7044 6134 7046
rect 5826 7035 6134 7044
rect 5172 6928 5224 6934
rect 4724 6886 4844 6914
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3896 5658 3924 6394
rect 3988 5846 4016 6598
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 3896 5630 4016 5658
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3804 3738 3832 4694
rect 3896 4690 3924 5034
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3988 4622 4016 5630
rect 4172 5370 4200 6802
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4264 5370 4292 6598
rect 4356 6458 4384 6886
rect 4469 6556 4777 6565
rect 4469 6554 4475 6556
rect 4531 6554 4555 6556
rect 4611 6554 4635 6556
rect 4691 6554 4715 6556
rect 4771 6554 4777 6556
rect 4531 6502 4533 6554
rect 4713 6502 4715 6554
rect 4469 6500 4475 6502
rect 4531 6500 4555 6502
rect 4611 6500 4635 6502
rect 4691 6500 4715 6502
rect 4771 6500 4777 6502
rect 4469 6491 4777 6500
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4816 5778 4844 6886
rect 6932 6882 6960 7890
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7024 7410 7052 7686
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7116 7342 7144 7822
rect 8036 7750 8064 7958
rect 8128 7818 8156 8366
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7183 7644 7491 7653
rect 7183 7642 7189 7644
rect 7245 7642 7269 7644
rect 7325 7642 7349 7644
rect 7405 7642 7429 7644
rect 7485 7642 7491 7644
rect 7245 7590 7247 7642
rect 7427 7590 7429 7642
rect 7183 7588 7189 7590
rect 7245 7588 7269 7590
rect 7325 7588 7349 7590
rect 7405 7588 7429 7590
rect 7485 7588 7491 7590
rect 7183 7579 7491 7588
rect 8036 7342 8064 7686
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7116 6914 7144 7278
rect 7760 7002 7788 7278
rect 8128 7206 8156 7754
rect 8312 7342 8340 8230
rect 8540 8188 8848 8197
rect 8540 8186 8546 8188
rect 8602 8186 8626 8188
rect 8682 8186 8706 8188
rect 8762 8186 8786 8188
rect 8842 8186 8848 8188
rect 8602 8134 8604 8186
rect 8784 8134 8786 8186
rect 8540 8132 8546 8134
rect 8602 8132 8626 8134
rect 8682 8132 8706 8134
rect 8762 8132 8786 8134
rect 8842 8132 8848 8134
rect 8540 8123 8848 8132
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 5172 6870 5224 6876
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4908 6390 4936 6802
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 4908 5914 4936 6326
rect 5184 6254 5212 6870
rect 6840 6854 6960 6882
rect 7024 6886 7144 6914
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 5276 6458 5304 6734
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5368 6338 5396 6394
rect 5276 6322 5396 6338
rect 5264 6316 5396 6322
rect 5316 6310 5396 6316
rect 5264 6258 5316 6264
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5184 5914 5212 6190
rect 5826 6012 6134 6021
rect 5826 6010 5832 6012
rect 5888 6010 5912 6012
rect 5968 6010 5992 6012
rect 6048 6010 6072 6012
rect 6128 6010 6134 6012
rect 5888 5958 5890 6010
rect 6070 5958 6072 6010
rect 5826 5956 5832 5958
rect 5888 5956 5912 5958
rect 5968 5956 5992 5958
rect 6048 5956 6072 5958
rect 6128 5956 6134 5958
rect 5826 5947 6134 5956
rect 6564 5914 6592 6734
rect 6840 6458 6868 6854
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4469 5468 4777 5477
rect 4469 5466 4475 5468
rect 4531 5466 4555 5468
rect 4611 5466 4635 5468
rect 4691 5466 4715 5468
rect 4771 5466 4777 5468
rect 4531 5414 4533 5466
rect 4713 5414 4715 5466
rect 4469 5412 4475 5414
rect 4531 5412 4555 5414
rect 4611 5412 4635 5414
rect 4691 5412 4715 5414
rect 4771 5412 4777 5414
rect 4469 5403 4777 5412
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3988 4146 4016 4558
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3804 3058 3832 3674
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3988 2922 4016 4082
rect 4264 4078 4292 5306
rect 4712 5092 4764 5098
rect 4816 5080 4844 5714
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 4764 5052 4844 5080
rect 4712 5034 4764 5040
rect 5000 5030 5028 5510
rect 6368 5296 6420 5302
rect 6368 5238 6420 5244
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 5826 4924 6134 4933
rect 5826 4922 5832 4924
rect 5888 4922 5912 4924
rect 5968 4922 5992 4924
rect 6048 4922 6072 4924
rect 6128 4922 6134 4924
rect 5888 4870 5890 4922
rect 6070 4870 6072 4922
rect 5826 4868 5832 4870
rect 5888 4868 5912 4870
rect 5968 4868 5992 4870
rect 6048 4868 6072 4870
rect 6128 4868 6134 4870
rect 5826 4859 6134 4868
rect 6196 4826 6224 5034
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6380 4690 6408 5238
rect 6932 5098 6960 6190
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 4690 6868 4966
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 4469 4380 4777 4389
rect 4469 4378 4475 4380
rect 4531 4378 4555 4380
rect 4611 4378 4635 4380
rect 4691 4378 4715 4380
rect 4771 4378 4777 4380
rect 4531 4326 4533 4378
rect 4713 4326 4715 4378
rect 4469 4324 4475 4326
rect 4531 4324 4555 4326
rect 4611 4324 4635 4326
rect 4691 4324 4715 4326
rect 4771 4324 4777 4326
rect 4469 4315 4777 4324
rect 6380 4078 6408 4626
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4469 3292 4777 3301
rect 4469 3290 4475 3292
rect 4531 3290 4555 3292
rect 4611 3290 4635 3292
rect 4691 3290 4715 3292
rect 4771 3290 4777 3292
rect 4531 3238 4533 3290
rect 4713 3238 4715 3290
rect 4469 3236 4475 3238
rect 4531 3236 4555 3238
rect 4611 3236 4635 3238
rect 4691 3236 4715 3238
rect 4771 3236 4777 3238
rect 4469 3227 4777 3236
rect 4816 2922 4844 3878
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4908 3058 4936 3334
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 3976 2916 4028 2922
rect 3976 2858 4028 2864
rect 4804 2916 4856 2922
rect 4804 2858 4856 2864
rect 4469 2204 4777 2213
rect 4469 2202 4475 2204
rect 4531 2202 4555 2204
rect 4611 2202 4635 2204
rect 4691 2202 4715 2204
rect 4771 2202 4777 2204
rect 4531 2150 4533 2202
rect 4713 2150 4715 2202
rect 4469 2148 4475 2150
rect 4531 2148 4555 2150
rect 4611 2148 4635 2150
rect 4691 2148 4715 2150
rect 4771 2148 4777 2150
rect 4469 2139 4777 2148
rect 1492 2100 1544 2106
rect 1492 2042 1544 2048
rect 3700 2100 3752 2106
rect 3700 2042 3752 2048
rect 4816 1970 4844 2858
rect 5644 2514 5672 4014
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 5826 3836 6134 3845
rect 5826 3834 5832 3836
rect 5888 3834 5912 3836
rect 5968 3834 5992 3836
rect 6048 3834 6072 3836
rect 6128 3834 6134 3836
rect 5888 3782 5890 3834
rect 6070 3782 6072 3834
rect 5826 3780 5832 3782
rect 5888 3780 5912 3782
rect 5968 3780 5992 3782
rect 6048 3780 6072 3782
rect 6128 3780 6134 3782
rect 5826 3771 6134 3780
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5092 2106 5120 2450
rect 5736 2446 5764 3538
rect 6196 2990 6224 3878
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 5826 2748 6134 2757
rect 5826 2746 5832 2748
rect 5888 2746 5912 2748
rect 5968 2746 5992 2748
rect 6048 2746 6072 2748
rect 6128 2746 6134 2748
rect 5888 2694 5890 2746
rect 6070 2694 6072 2746
rect 5826 2692 5832 2694
rect 5888 2692 5912 2694
rect 5968 2692 5992 2694
rect 6048 2692 6072 2694
rect 6128 2692 6134 2694
rect 5826 2683 6134 2692
rect 6380 2650 6408 4014
rect 6932 3942 6960 5034
rect 7024 5030 7052 6886
rect 7116 6730 7144 6886
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7183 6556 7491 6565
rect 7183 6554 7189 6556
rect 7245 6554 7269 6556
rect 7325 6554 7349 6556
rect 7405 6554 7429 6556
rect 7485 6554 7491 6556
rect 7245 6502 7247 6554
rect 7427 6502 7429 6554
rect 7183 6500 7189 6502
rect 7245 6500 7269 6502
rect 7325 6500 7349 6502
rect 7405 6500 7429 6502
rect 7485 6500 7491 6502
rect 7183 6491 7491 6500
rect 7668 6458 7696 6802
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7564 6180 7616 6186
rect 7564 6122 7616 6128
rect 7576 6089 7604 6122
rect 7562 6080 7618 6089
rect 7562 6015 7618 6024
rect 7760 5914 7788 6938
rect 8024 6928 8076 6934
rect 8220 6914 8248 7142
rect 8300 6928 8352 6934
rect 8220 6886 8300 6914
rect 8024 6870 8076 6876
rect 8300 6870 8352 6876
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7183 5468 7491 5477
rect 7183 5466 7189 5468
rect 7245 5466 7269 5468
rect 7325 5466 7349 5468
rect 7405 5466 7429 5468
rect 7485 5466 7491 5468
rect 7245 5414 7247 5466
rect 7427 5414 7429 5466
rect 7183 5412 7189 5414
rect 7245 5412 7269 5414
rect 7325 5412 7349 5414
rect 7405 5412 7429 5414
rect 7485 5412 7491 5414
rect 7183 5403 7491 5412
rect 7668 5234 7696 5714
rect 7852 5710 7880 6054
rect 8036 5914 8064 6870
rect 8404 6662 8432 7414
rect 8588 7342 8616 7686
rect 8956 7546 8984 8298
rect 9048 7954 9076 8366
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8540 7100 8848 7109
rect 8540 7098 8546 7100
rect 8602 7098 8626 7100
rect 8682 7098 8706 7100
rect 8762 7098 8786 7100
rect 8842 7098 8848 7100
rect 8602 7046 8604 7098
rect 8784 7046 8786 7098
rect 8540 7044 8546 7046
rect 8602 7044 8626 7046
rect 8682 7044 8706 7046
rect 8762 7044 8786 7046
rect 8842 7044 8848 7046
rect 8540 7035 8848 7044
rect 9048 6866 9076 7686
rect 9140 7410 9168 8230
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9324 7546 9352 7890
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9140 7002 9168 7346
rect 9416 7342 9444 8570
rect 11254 8188 11562 8197
rect 11254 8186 11260 8188
rect 11316 8186 11340 8188
rect 11396 8186 11420 8188
rect 11476 8186 11500 8188
rect 11556 8186 11562 8188
rect 11316 8134 11318 8186
rect 11498 8134 11500 8186
rect 11254 8132 11260 8134
rect 11316 8132 11340 8134
rect 11396 8132 11420 8134
rect 11476 8132 11500 8134
rect 11556 8132 11562 8134
rect 11254 8123 11562 8132
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 9897 7644 10205 7653
rect 9897 7642 9903 7644
rect 9959 7642 9983 7644
rect 10039 7642 10063 7644
rect 10119 7642 10143 7644
rect 10199 7642 10205 7644
rect 9959 7590 9961 7642
rect 10141 7590 10143 7642
rect 9897 7588 9903 7590
rect 9959 7588 9983 7590
rect 10039 7588 10063 7590
rect 10119 7588 10143 7590
rect 10199 7588 10205 7590
rect 9897 7579 10205 7588
rect 10612 7410 10640 7686
rect 11058 7440 11114 7449
rect 10600 7404 10652 7410
rect 11058 7375 11114 7384
rect 10600 7346 10652 7352
rect 11072 7342 11100 7375
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 10888 6866 10916 7142
rect 11254 7100 11562 7109
rect 11254 7098 11260 7100
rect 11316 7098 11340 7100
rect 11396 7098 11420 7100
rect 11476 7098 11500 7100
rect 11556 7098 11562 7100
rect 11316 7046 11318 7098
rect 11498 7046 11500 7098
rect 11254 7044 11260 7046
rect 11316 7044 11340 7046
rect 11396 7044 11420 7046
rect 11476 7044 11500 7046
rect 11556 7044 11562 7046
rect 11254 7035 11562 7044
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 8220 5778 8248 6598
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8312 5914 8340 6190
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8404 5794 8432 6598
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8540 6012 8848 6021
rect 8540 6010 8546 6012
rect 8602 6010 8626 6012
rect 8682 6010 8706 6012
rect 8762 6010 8786 6012
rect 8842 6010 8848 6012
rect 8602 5958 8604 6010
rect 8784 5958 8786 6010
rect 8540 5956 8546 5958
rect 8602 5956 8626 5958
rect 8682 5956 8706 5958
rect 8762 5956 8786 5958
rect 8842 5956 8848 5958
rect 8540 5947 8848 5956
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8312 5766 8432 5794
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7024 4758 7052 4966
rect 7484 4826 7512 4966
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 7183 4380 7491 4389
rect 7183 4378 7189 4380
rect 7245 4378 7269 4380
rect 7325 4378 7349 4380
rect 7405 4378 7429 4380
rect 7485 4378 7491 4380
rect 7245 4326 7247 4378
rect 7427 4326 7429 4378
rect 7183 4324 7189 4326
rect 7245 4324 7269 4326
rect 7325 4324 7349 4326
rect 7405 4324 7429 4326
rect 7485 4324 7491 4326
rect 7183 4315 7491 4324
rect 7668 4214 7696 5170
rect 7760 5166 7788 5646
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7760 4282 7788 5102
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7656 4208 7708 4214
rect 7656 4150 7708 4156
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 7760 3602 7788 4014
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 6656 2990 6684 3538
rect 7183 3292 7491 3301
rect 7183 3290 7189 3292
rect 7245 3290 7269 3292
rect 7325 3290 7349 3292
rect 7405 3290 7429 3292
rect 7485 3290 7491 3292
rect 7245 3238 7247 3290
rect 7427 3238 7429 3290
rect 7183 3236 7189 3238
rect 7245 3236 7269 3238
rect 7325 3236 7349 3238
rect 7405 3236 7429 3238
rect 7485 3236 7491 3238
rect 7183 3227 7491 3236
rect 7760 3194 7788 3538
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 7852 3074 7880 5646
rect 8312 5166 8340 5766
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5234 8524 5510
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8128 4826 8156 5034
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 7944 3602 7972 4014
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7944 3398 7972 3538
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 8036 3346 8064 3878
rect 8128 3738 8156 4014
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8220 3602 8248 4014
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8312 3534 8340 4082
rect 8404 3670 8432 5102
rect 8540 4924 8848 4933
rect 8540 4922 8546 4924
rect 8602 4922 8626 4924
rect 8682 4922 8706 4924
rect 8762 4922 8786 4924
rect 8842 4922 8848 4924
rect 8602 4870 8604 4922
rect 8784 4870 8786 4922
rect 8540 4868 8546 4870
rect 8602 4868 8626 4870
rect 8682 4868 8706 4870
rect 8762 4868 8786 4870
rect 8842 4868 8848 4870
rect 8540 4859 8848 4868
rect 8956 4146 8984 6190
rect 9600 5778 9628 6666
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6186 9720 6598
rect 9784 6440 9812 6802
rect 9897 6556 10205 6565
rect 9897 6554 9903 6556
rect 9959 6554 9983 6556
rect 10039 6554 10063 6556
rect 10119 6554 10143 6556
rect 10199 6554 10205 6556
rect 9959 6502 9961 6554
rect 10141 6502 10143 6554
rect 9897 6500 9903 6502
rect 9959 6500 9983 6502
rect 10039 6500 10063 6502
rect 10119 6500 10143 6502
rect 10199 6500 10205 6502
rect 9897 6491 10205 6500
rect 9784 6412 9904 6440
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 9140 4078 9168 4626
rect 9508 4162 9536 5306
rect 9600 5098 9628 5510
rect 9588 5092 9640 5098
rect 9588 5034 9640 5040
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9416 4146 9628 4162
rect 9416 4140 9640 4146
rect 9416 4134 9588 4140
rect 8760 4072 8812 4078
rect 9036 4072 9088 4078
rect 8812 4020 8984 4026
rect 8760 4014 8984 4020
rect 9036 4014 9088 4020
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 8772 3998 8984 4014
rect 8540 3836 8848 3845
rect 8540 3834 8546 3836
rect 8602 3834 8626 3836
rect 8682 3834 8706 3836
rect 8762 3834 8786 3836
rect 8842 3834 8848 3836
rect 8602 3782 8604 3834
rect 8784 3782 8786 3834
rect 8540 3780 8546 3782
rect 8602 3780 8626 3782
rect 8682 3780 8706 3782
rect 8762 3780 8786 3782
rect 8842 3780 8848 3782
rect 8540 3771 8848 3780
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8036 3318 8248 3346
rect 8220 3126 8248 3318
rect 8496 3194 8524 3538
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 7760 3046 7880 3074
rect 8208 3120 8260 3126
rect 8588 3074 8616 3470
rect 8208 3062 8260 3068
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 7760 2650 7788 3046
rect 8220 2774 8248 3062
rect 8496 3058 8616 3074
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 8484 3052 8616 3058
rect 8536 3046 8616 3052
rect 8484 2994 8536 3000
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8588 2938 8616 3046
rect 8864 2990 8892 3062
rect 8852 2984 8904 2990
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8128 2746 8248 2774
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 5080 2100 5132 2106
rect 5080 2042 5132 2048
rect 5368 1970 5396 2246
rect 6012 1970 6040 2450
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 4804 1964 4856 1970
rect 4804 1906 4856 1912
rect 5356 1964 5408 1970
rect 5356 1906 5408 1912
rect 6000 1964 6052 1970
rect 6000 1906 6052 1912
rect 2688 1828 2740 1834
rect 2688 1770 2740 1776
rect 3516 1828 3568 1834
rect 3516 1770 3568 1776
rect 2700 1562 2728 1770
rect 3112 1660 3420 1669
rect 3112 1658 3118 1660
rect 3174 1658 3198 1660
rect 3254 1658 3278 1660
rect 3334 1658 3358 1660
rect 3414 1658 3420 1660
rect 3174 1606 3176 1658
rect 3356 1606 3358 1658
rect 3112 1604 3118 1606
rect 3174 1604 3198 1606
rect 3254 1604 3278 1606
rect 3334 1604 3358 1606
rect 3414 1604 3420 1606
rect 3112 1595 3420 1604
rect 3528 1562 3556 1770
rect 2688 1556 2740 1562
rect 2688 1498 2740 1504
rect 3516 1556 3568 1562
rect 3516 1498 3568 1504
rect 1400 1420 1452 1426
rect 1400 1362 1452 1368
rect 1412 1018 1440 1362
rect 4816 1358 4844 1906
rect 6104 1834 6132 2246
rect 7183 2204 7491 2213
rect 7183 2202 7189 2204
rect 7245 2202 7269 2204
rect 7325 2202 7349 2204
rect 7405 2202 7429 2204
rect 7485 2202 7491 2204
rect 7245 2150 7247 2202
rect 7427 2150 7429 2202
rect 7183 2148 7189 2150
rect 7245 2148 7269 2150
rect 7325 2148 7349 2150
rect 7405 2148 7429 2150
rect 7485 2148 7491 2150
rect 7183 2139 7491 2148
rect 7760 1902 7788 2586
rect 8128 2394 8156 2746
rect 8312 2582 8340 2858
rect 8404 2582 8432 2926
rect 8588 2910 8800 2938
rect 8852 2926 8904 2932
rect 8772 2854 8800 2910
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8540 2748 8848 2757
rect 8540 2746 8546 2748
rect 8602 2746 8626 2748
rect 8682 2746 8706 2748
rect 8762 2746 8786 2748
rect 8842 2746 8848 2748
rect 8602 2694 8604 2746
rect 8784 2694 8786 2746
rect 8540 2692 8546 2694
rect 8602 2692 8626 2694
rect 8682 2692 8706 2694
rect 8762 2692 8786 2694
rect 8842 2692 8848 2694
rect 8540 2683 8848 2692
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8392 2576 8444 2582
rect 8392 2518 8444 2524
rect 8300 2440 8352 2446
rect 8128 2388 8300 2394
rect 8956 2394 8984 3998
rect 9048 3738 9076 4014
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 9048 3602 9076 3674
rect 9324 3602 9352 4014
rect 9036 3596 9088 3602
rect 9312 3596 9364 3602
rect 9036 3538 9088 3544
rect 9232 3556 9312 3584
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9140 3058 9168 3470
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9048 2650 9076 2926
rect 9140 2854 9168 2994
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9232 2530 9260 3556
rect 9312 3538 9364 3544
rect 9416 3398 9444 4134
rect 9588 4082 9640 4088
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9416 3194 9444 3334
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9416 2938 9444 3130
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9600 3074 9628 3538
rect 9692 3194 9720 4558
rect 9784 4282 9812 6054
rect 9876 5846 9904 6412
rect 10428 6254 10456 6802
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9897 5468 10205 5477
rect 9897 5466 9903 5468
rect 9959 5466 9983 5468
rect 10039 5466 10063 5468
rect 10119 5466 10143 5468
rect 10199 5466 10205 5468
rect 9959 5414 9961 5466
rect 10141 5414 10143 5466
rect 9897 5412 9903 5414
rect 9959 5412 9983 5414
rect 10039 5412 10063 5414
rect 10119 5412 10143 5414
rect 10199 5412 10205 5414
rect 9897 5403 10205 5412
rect 10428 5166 10456 6190
rect 11254 6012 11562 6021
rect 11254 6010 11260 6012
rect 11316 6010 11340 6012
rect 11396 6010 11420 6012
rect 11476 6010 11500 6012
rect 11556 6010 11562 6012
rect 11316 5958 11318 6010
rect 11498 5958 11500 6010
rect 11254 5956 11260 5958
rect 11316 5956 11340 5958
rect 11396 5956 11420 5958
rect 11476 5956 11500 5958
rect 11556 5956 11562 5958
rect 11254 5947 11562 5956
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10244 4758 10272 4966
rect 11254 4924 11562 4933
rect 11254 4922 11260 4924
rect 11316 4922 11340 4924
rect 11396 4922 11420 4924
rect 11476 4922 11500 4924
rect 11556 4922 11562 4924
rect 11316 4870 11318 4922
rect 11498 4870 11500 4922
rect 11254 4868 11260 4870
rect 11316 4868 11340 4870
rect 11396 4868 11420 4870
rect 11476 4868 11500 4870
rect 11556 4868 11562 4870
rect 11254 4859 11562 4868
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 9897 4380 10205 4389
rect 9897 4378 9903 4380
rect 9959 4378 9983 4380
rect 10039 4378 10063 4380
rect 10119 4378 10143 4380
rect 10199 4378 10205 4380
rect 9959 4326 9961 4378
rect 10141 4326 10143 4378
rect 9897 4324 9903 4326
rect 9959 4324 9983 4326
rect 10039 4324 10063 4326
rect 10119 4324 10143 4326
rect 10199 4324 10205 4326
rect 9897 4315 10205 4324
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9784 4078 9812 4218
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 10244 3602 10272 4694
rect 11254 3836 11562 3845
rect 11254 3834 11260 3836
rect 11316 3834 11340 3836
rect 11396 3834 11420 3836
rect 11476 3834 11500 3836
rect 11556 3834 11562 3836
rect 11316 3782 11318 3834
rect 11498 3782 11500 3834
rect 11254 3780 11260 3782
rect 11316 3780 11340 3782
rect 11396 3780 11420 3782
rect 11476 3780 11500 3782
rect 11556 3780 11562 3782
rect 11254 3771 11562 3780
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 9897 3292 10205 3301
rect 9897 3290 9903 3292
rect 9959 3290 9983 3292
rect 10039 3290 10063 3292
rect 10119 3290 10143 3292
rect 10199 3290 10205 3292
rect 9959 3238 9961 3290
rect 10141 3238 10143 3290
rect 9897 3236 9903 3238
rect 9959 3236 9983 3238
rect 10039 3236 10063 3238
rect 10119 3236 10143 3238
rect 10199 3236 10205 3238
rect 9897 3227 10205 3236
rect 10428 3194 10456 3470
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 9876 3074 9904 3130
rect 9140 2514 9260 2530
rect 9128 2508 9260 2514
rect 9180 2502 9260 2508
rect 9324 2910 9444 2938
rect 9508 2938 9536 3062
rect 9600 3046 9904 3074
rect 9508 2922 9720 2938
rect 9508 2916 9732 2922
rect 9508 2910 9680 2916
rect 9128 2450 9180 2456
rect 8128 2382 8352 2388
rect 8128 2366 8340 2382
rect 7748 1896 7800 1902
rect 7748 1838 7800 1844
rect 6092 1828 6144 1834
rect 6092 1770 6144 1776
rect 7196 1760 7248 1766
rect 7196 1702 7248 1708
rect 5826 1660 6134 1669
rect 5826 1658 5832 1660
rect 5888 1658 5912 1660
rect 5968 1658 5992 1660
rect 6048 1658 6072 1660
rect 6128 1658 6134 1660
rect 5888 1606 5890 1658
rect 6070 1606 6072 1658
rect 5826 1604 5832 1606
rect 5888 1604 5912 1606
rect 5968 1604 5992 1606
rect 6048 1604 6072 1606
rect 6128 1604 6134 1606
rect 5826 1595 6134 1604
rect 7208 1494 7236 1702
rect 7760 1562 7788 1838
rect 7748 1556 7800 1562
rect 7748 1498 7800 1504
rect 7196 1488 7248 1494
rect 7196 1430 7248 1436
rect 8312 1426 8340 2366
rect 8864 2366 8984 2394
rect 8864 2310 8892 2366
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 8864 1902 8892 2246
rect 9232 2038 9260 2246
rect 9324 2106 9352 2910
rect 9680 2858 9732 2864
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9416 2310 9444 2790
rect 9508 2378 9536 2790
rect 9876 2650 9904 3046
rect 11254 2748 11562 2757
rect 11254 2746 11260 2748
rect 11316 2746 11340 2748
rect 11396 2746 11420 2748
rect 11476 2746 11500 2748
rect 11556 2746 11562 2748
rect 11316 2694 11318 2746
rect 11498 2694 11500 2746
rect 11254 2692 11260 2694
rect 11316 2692 11340 2694
rect 11396 2692 11420 2694
rect 11476 2692 11500 2694
rect 11556 2692 11562 2694
rect 11254 2683 11562 2692
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9496 2372 9548 2378
rect 9496 2314 9548 2320
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9897 2204 10205 2213
rect 9897 2202 9903 2204
rect 9959 2202 9983 2204
rect 10039 2202 10063 2204
rect 10119 2202 10143 2204
rect 10199 2202 10205 2204
rect 9959 2150 9961 2202
rect 10141 2150 10143 2202
rect 9897 2148 9903 2150
rect 9959 2148 9983 2150
rect 10039 2148 10063 2150
rect 10119 2148 10143 2150
rect 10199 2148 10205 2150
rect 9897 2139 10205 2148
rect 9312 2100 9364 2106
rect 9312 2042 9364 2048
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 8852 1896 8904 1902
rect 8852 1838 8904 1844
rect 8392 1760 8444 1766
rect 8392 1702 8444 1708
rect 5540 1420 5592 1426
rect 5540 1362 5592 1368
rect 8300 1420 8352 1426
rect 8300 1362 8352 1368
rect 4068 1352 4120 1358
rect 4068 1294 4120 1300
rect 4804 1352 4856 1358
rect 4804 1294 4856 1300
rect 3332 1216 3384 1222
rect 3332 1158 3384 1164
rect 1755 1116 2063 1125
rect 1755 1114 1761 1116
rect 1817 1114 1841 1116
rect 1897 1114 1921 1116
rect 1977 1114 2001 1116
rect 2057 1114 2063 1116
rect 1817 1062 1819 1114
rect 1999 1062 2001 1114
rect 1755 1060 1761 1062
rect 1817 1060 1841 1062
rect 1897 1060 1921 1062
rect 1977 1060 2001 1062
rect 2057 1060 2063 1062
rect 1755 1051 2063 1060
rect 3344 1018 3372 1158
rect 1400 1012 1452 1018
rect 1400 954 1452 960
rect 3332 1012 3384 1018
rect 3332 954 3384 960
rect 4080 950 4108 1294
rect 4469 1116 4777 1125
rect 4469 1114 4475 1116
rect 4531 1114 4555 1116
rect 4611 1114 4635 1116
rect 4691 1114 4715 1116
rect 4771 1114 4777 1116
rect 4531 1062 4533 1114
rect 4713 1062 4715 1114
rect 4469 1060 4475 1062
rect 4531 1060 4555 1062
rect 4611 1060 4635 1062
rect 4691 1060 4715 1062
rect 4771 1060 4777 1062
rect 4469 1051 4777 1060
rect 5552 1018 5580 1362
rect 8404 1358 8432 1702
rect 8540 1660 8848 1669
rect 8540 1658 8546 1660
rect 8602 1658 8626 1660
rect 8682 1658 8706 1660
rect 8762 1658 8786 1660
rect 8842 1658 8848 1660
rect 8602 1606 8604 1658
rect 8784 1606 8786 1658
rect 8540 1604 8546 1606
rect 8602 1604 8626 1606
rect 8682 1604 8706 1606
rect 8762 1604 8786 1606
rect 8842 1604 8848 1606
rect 8540 1595 8848 1604
rect 11254 1660 11562 1669
rect 11254 1658 11260 1660
rect 11316 1658 11340 1660
rect 11396 1658 11420 1660
rect 11476 1658 11500 1660
rect 11556 1658 11562 1660
rect 11316 1606 11318 1658
rect 11498 1606 11500 1658
rect 11254 1604 11260 1606
rect 11316 1604 11340 1606
rect 11396 1604 11420 1606
rect 11476 1604 11500 1606
rect 11556 1604 11562 1606
rect 11254 1595 11562 1604
rect 10692 1420 10744 1426
rect 10692 1362 10744 1368
rect 8392 1352 8444 1358
rect 8392 1294 8444 1300
rect 7183 1116 7491 1125
rect 7183 1114 7189 1116
rect 7245 1114 7269 1116
rect 7325 1114 7349 1116
rect 7405 1114 7429 1116
rect 7485 1114 7491 1116
rect 7245 1062 7247 1114
rect 7427 1062 7429 1114
rect 7183 1060 7189 1062
rect 7245 1060 7269 1062
rect 7325 1060 7349 1062
rect 7405 1060 7429 1062
rect 7485 1060 7491 1062
rect 7183 1051 7491 1060
rect 9897 1116 10205 1125
rect 9897 1114 9903 1116
rect 9959 1114 9983 1116
rect 10039 1114 10063 1116
rect 10119 1114 10143 1116
rect 10199 1114 10205 1116
rect 9959 1062 9961 1114
rect 10141 1062 10143 1114
rect 9897 1060 9903 1062
rect 9959 1060 9983 1062
rect 10039 1060 10063 1062
rect 10119 1060 10143 1062
rect 10199 1060 10205 1062
rect 9897 1051 10205 1060
rect 5540 1012 5592 1018
rect 5540 954 5592 960
rect 4068 944 4120 950
rect 4068 886 4120 892
rect 1124 808 1176 814
rect 1124 750 1176 756
rect 3516 808 3568 814
rect 3516 750 3568 756
rect 6184 808 6236 814
rect 6184 750 6236 756
rect 8300 808 8352 814
rect 8300 750 8352 756
rect 1136 400 1164 750
rect 3112 572 3420 581
rect 3112 570 3118 572
rect 3174 570 3198 572
rect 3254 570 3278 572
rect 3334 570 3358 572
rect 3414 570 3420 572
rect 3174 518 3176 570
rect 3356 518 3358 570
rect 3112 516 3118 518
rect 3174 516 3198 518
rect 3254 516 3278 518
rect 3334 516 3358 518
rect 3414 516 3420 518
rect 3112 507 3420 516
rect 3528 400 3556 750
rect 5826 572 6134 581
rect 5826 570 5832 572
rect 5888 570 5912 572
rect 5968 570 5992 572
rect 6048 570 6072 572
rect 6128 570 6134 572
rect 5888 518 5890 570
rect 6070 518 6072 570
rect 5826 516 5832 518
rect 5888 516 5912 518
rect 5968 516 5992 518
rect 6048 516 6072 518
rect 6128 516 6134 518
rect 5826 507 6134 516
rect 6196 456 6224 750
rect 5920 428 6224 456
rect 5920 400 5948 428
rect 8312 400 8340 750
rect 8540 572 8848 581
rect 8540 570 8546 572
rect 8602 570 8626 572
rect 8682 570 8706 572
rect 8762 570 8786 572
rect 8842 570 8848 572
rect 8602 518 8604 570
rect 8784 518 8786 570
rect 8540 516 8546 518
rect 8602 516 8626 518
rect 8682 516 8706 518
rect 8762 516 8786 518
rect 8842 516 8848 518
rect 8540 507 8848 516
rect 10704 400 10732 1362
rect 11254 572 11562 581
rect 11254 570 11260 572
rect 11316 570 11340 572
rect 11396 570 11420 572
rect 11476 570 11500 572
rect 11556 570 11562 572
rect 11316 518 11318 570
rect 11498 518 11500 570
rect 11254 516 11260 518
rect 11316 516 11340 518
rect 11396 516 11420 518
rect 11476 516 11500 518
rect 11556 516 11562 518
rect 11254 507 11562 516
rect 1122 0 1178 400
rect 3514 0 3570 400
rect 5906 0 5962 400
rect 8298 0 8354 400
rect 10690 0 10746 400
<< via2 >>
rect 3118 9274 3174 9276
rect 3198 9274 3254 9276
rect 3278 9274 3334 9276
rect 3358 9274 3414 9276
rect 3118 9222 3164 9274
rect 3164 9222 3174 9274
rect 3198 9222 3228 9274
rect 3228 9222 3240 9274
rect 3240 9222 3254 9274
rect 3278 9222 3292 9274
rect 3292 9222 3304 9274
rect 3304 9222 3334 9274
rect 3358 9222 3368 9274
rect 3368 9222 3414 9274
rect 3118 9220 3174 9222
rect 3198 9220 3254 9222
rect 3278 9220 3334 9222
rect 3358 9220 3414 9222
rect 1761 8730 1817 8732
rect 1841 8730 1897 8732
rect 1921 8730 1977 8732
rect 2001 8730 2057 8732
rect 1761 8678 1807 8730
rect 1807 8678 1817 8730
rect 1841 8678 1871 8730
rect 1871 8678 1883 8730
rect 1883 8678 1897 8730
rect 1921 8678 1935 8730
rect 1935 8678 1947 8730
rect 1947 8678 1977 8730
rect 2001 8678 2011 8730
rect 2011 8678 2057 8730
rect 1761 8676 1817 8678
rect 1841 8676 1897 8678
rect 1921 8676 1977 8678
rect 2001 8676 2057 8678
rect 3118 8186 3174 8188
rect 3198 8186 3254 8188
rect 3278 8186 3334 8188
rect 3358 8186 3414 8188
rect 3118 8134 3164 8186
rect 3164 8134 3174 8186
rect 3198 8134 3228 8186
rect 3228 8134 3240 8186
rect 3240 8134 3254 8186
rect 3278 8134 3292 8186
rect 3292 8134 3304 8186
rect 3304 8134 3334 8186
rect 3358 8134 3368 8186
rect 3368 8134 3414 8186
rect 3118 8132 3174 8134
rect 3198 8132 3254 8134
rect 3278 8132 3334 8134
rect 3358 8132 3414 8134
rect 1761 7642 1817 7644
rect 1841 7642 1897 7644
rect 1921 7642 1977 7644
rect 2001 7642 2057 7644
rect 1761 7590 1807 7642
rect 1807 7590 1817 7642
rect 1841 7590 1871 7642
rect 1871 7590 1883 7642
rect 1883 7590 1897 7642
rect 1921 7590 1935 7642
rect 1935 7590 1947 7642
rect 1947 7590 1977 7642
rect 2001 7590 2011 7642
rect 2011 7590 2057 7642
rect 1761 7588 1817 7590
rect 1841 7588 1897 7590
rect 1921 7588 1977 7590
rect 2001 7588 2057 7590
rect 3118 7098 3174 7100
rect 3198 7098 3254 7100
rect 3278 7098 3334 7100
rect 3358 7098 3414 7100
rect 3118 7046 3164 7098
rect 3164 7046 3174 7098
rect 3198 7046 3228 7098
rect 3228 7046 3240 7098
rect 3240 7046 3254 7098
rect 3278 7046 3292 7098
rect 3292 7046 3304 7098
rect 3304 7046 3334 7098
rect 3358 7046 3368 7098
rect 3368 7046 3414 7098
rect 3118 7044 3174 7046
rect 3198 7044 3254 7046
rect 3278 7044 3334 7046
rect 3358 7044 3414 7046
rect 1761 6554 1817 6556
rect 1841 6554 1897 6556
rect 1921 6554 1977 6556
rect 2001 6554 2057 6556
rect 1761 6502 1807 6554
rect 1807 6502 1817 6554
rect 1841 6502 1871 6554
rect 1871 6502 1883 6554
rect 1883 6502 1897 6554
rect 1921 6502 1935 6554
rect 1935 6502 1947 6554
rect 1947 6502 1977 6554
rect 2001 6502 2011 6554
rect 2011 6502 2057 6554
rect 1761 6500 1817 6502
rect 1841 6500 1897 6502
rect 1921 6500 1977 6502
rect 2001 6500 2057 6502
rect 1761 5466 1817 5468
rect 1841 5466 1897 5468
rect 1921 5466 1977 5468
rect 2001 5466 2057 5468
rect 1761 5414 1807 5466
rect 1807 5414 1817 5466
rect 1841 5414 1871 5466
rect 1871 5414 1883 5466
rect 1883 5414 1897 5466
rect 1921 5414 1935 5466
rect 1935 5414 1947 5466
rect 1947 5414 1977 5466
rect 2001 5414 2011 5466
rect 2011 5414 2057 5466
rect 1761 5412 1817 5414
rect 1841 5412 1897 5414
rect 1921 5412 1977 5414
rect 2001 5412 2057 5414
rect 3118 6010 3174 6012
rect 3198 6010 3254 6012
rect 3278 6010 3334 6012
rect 3358 6010 3414 6012
rect 3118 5958 3164 6010
rect 3164 5958 3174 6010
rect 3198 5958 3228 6010
rect 3228 5958 3240 6010
rect 3240 5958 3254 6010
rect 3278 5958 3292 6010
rect 3292 5958 3304 6010
rect 3304 5958 3334 6010
rect 3358 5958 3368 6010
rect 3368 5958 3414 6010
rect 3118 5956 3174 5958
rect 3198 5956 3254 5958
rect 3278 5956 3334 5958
rect 3358 5956 3414 5958
rect 1761 4378 1817 4380
rect 1841 4378 1897 4380
rect 1921 4378 1977 4380
rect 2001 4378 2057 4380
rect 1761 4326 1807 4378
rect 1807 4326 1817 4378
rect 1841 4326 1871 4378
rect 1871 4326 1883 4378
rect 1883 4326 1897 4378
rect 1921 4326 1935 4378
rect 1935 4326 1947 4378
rect 1947 4326 1977 4378
rect 2001 4326 2011 4378
rect 2011 4326 2057 4378
rect 1761 4324 1817 4326
rect 1841 4324 1897 4326
rect 1921 4324 1977 4326
rect 2001 4324 2057 4326
rect 3118 4922 3174 4924
rect 3198 4922 3254 4924
rect 3278 4922 3334 4924
rect 3358 4922 3414 4924
rect 3118 4870 3164 4922
rect 3164 4870 3174 4922
rect 3198 4870 3228 4922
rect 3228 4870 3240 4922
rect 3240 4870 3254 4922
rect 3278 4870 3292 4922
rect 3292 4870 3304 4922
rect 3304 4870 3334 4922
rect 3358 4870 3368 4922
rect 3368 4870 3414 4922
rect 3118 4868 3174 4870
rect 3198 4868 3254 4870
rect 3278 4868 3334 4870
rect 3358 4868 3414 4870
rect 3118 3834 3174 3836
rect 3198 3834 3254 3836
rect 3278 3834 3334 3836
rect 3358 3834 3414 3836
rect 3118 3782 3164 3834
rect 3164 3782 3174 3834
rect 3198 3782 3228 3834
rect 3228 3782 3240 3834
rect 3240 3782 3254 3834
rect 3278 3782 3292 3834
rect 3292 3782 3304 3834
rect 3304 3782 3334 3834
rect 3358 3782 3368 3834
rect 3368 3782 3414 3834
rect 3118 3780 3174 3782
rect 3198 3780 3254 3782
rect 3278 3780 3334 3782
rect 3358 3780 3414 3782
rect 1761 3290 1817 3292
rect 1841 3290 1897 3292
rect 1921 3290 1977 3292
rect 2001 3290 2057 3292
rect 1761 3238 1807 3290
rect 1807 3238 1817 3290
rect 1841 3238 1871 3290
rect 1871 3238 1883 3290
rect 1883 3238 1897 3290
rect 1921 3238 1935 3290
rect 1935 3238 1947 3290
rect 1947 3238 1977 3290
rect 2001 3238 2011 3290
rect 2011 3238 2057 3290
rect 1761 3236 1817 3238
rect 1841 3236 1897 3238
rect 1921 3236 1977 3238
rect 2001 3236 2057 3238
rect 3118 2746 3174 2748
rect 3198 2746 3254 2748
rect 3278 2746 3334 2748
rect 3358 2746 3414 2748
rect 3118 2694 3164 2746
rect 3164 2694 3174 2746
rect 3198 2694 3228 2746
rect 3228 2694 3240 2746
rect 3240 2694 3254 2746
rect 3278 2694 3292 2746
rect 3292 2694 3304 2746
rect 3304 2694 3334 2746
rect 3358 2694 3368 2746
rect 3368 2694 3414 2746
rect 3118 2692 3174 2694
rect 3198 2692 3254 2694
rect 3278 2692 3334 2694
rect 3358 2692 3414 2694
rect 1761 2202 1817 2204
rect 1841 2202 1897 2204
rect 1921 2202 1977 2204
rect 2001 2202 2057 2204
rect 1761 2150 1807 2202
rect 1807 2150 1817 2202
rect 1841 2150 1871 2202
rect 1871 2150 1883 2202
rect 1883 2150 1897 2202
rect 1921 2150 1935 2202
rect 1935 2150 1947 2202
rect 1947 2150 1977 2202
rect 2001 2150 2011 2202
rect 2011 2150 2057 2202
rect 1761 2148 1817 2150
rect 1841 2148 1897 2150
rect 1921 2148 1977 2150
rect 2001 2148 2057 2150
rect 5832 9274 5888 9276
rect 5912 9274 5968 9276
rect 5992 9274 6048 9276
rect 6072 9274 6128 9276
rect 5832 9222 5878 9274
rect 5878 9222 5888 9274
rect 5912 9222 5942 9274
rect 5942 9222 5954 9274
rect 5954 9222 5968 9274
rect 5992 9222 6006 9274
rect 6006 9222 6018 9274
rect 6018 9222 6048 9274
rect 6072 9222 6082 9274
rect 6082 9222 6128 9274
rect 5832 9220 5888 9222
rect 5912 9220 5968 9222
rect 5992 9220 6048 9222
rect 6072 9220 6128 9222
rect 4475 8730 4531 8732
rect 4555 8730 4611 8732
rect 4635 8730 4691 8732
rect 4715 8730 4771 8732
rect 4475 8678 4521 8730
rect 4521 8678 4531 8730
rect 4555 8678 4585 8730
rect 4585 8678 4597 8730
rect 4597 8678 4611 8730
rect 4635 8678 4649 8730
rect 4649 8678 4661 8730
rect 4661 8678 4691 8730
rect 4715 8678 4725 8730
rect 4725 8678 4771 8730
rect 4475 8676 4531 8678
rect 4555 8676 4611 8678
rect 4635 8676 4691 8678
rect 4715 8676 4771 8678
rect 4475 7642 4531 7644
rect 4555 7642 4611 7644
rect 4635 7642 4691 7644
rect 4715 7642 4771 7644
rect 4475 7590 4521 7642
rect 4521 7590 4531 7642
rect 4555 7590 4585 7642
rect 4585 7590 4597 7642
rect 4597 7590 4611 7642
rect 4635 7590 4649 7642
rect 4649 7590 4661 7642
rect 4661 7590 4691 7642
rect 4715 7590 4725 7642
rect 4725 7590 4771 7642
rect 4475 7588 4531 7590
rect 4555 7588 4611 7590
rect 4635 7588 4691 7590
rect 4715 7588 4771 7590
rect 8546 9274 8602 9276
rect 8626 9274 8682 9276
rect 8706 9274 8762 9276
rect 8786 9274 8842 9276
rect 8546 9222 8592 9274
rect 8592 9222 8602 9274
rect 8626 9222 8656 9274
rect 8656 9222 8668 9274
rect 8668 9222 8682 9274
rect 8706 9222 8720 9274
rect 8720 9222 8732 9274
rect 8732 9222 8762 9274
rect 8786 9222 8796 9274
rect 8796 9222 8842 9274
rect 8546 9220 8602 9222
rect 8626 9220 8682 9222
rect 8706 9220 8762 9222
rect 8786 9220 8842 9222
rect 7189 8730 7245 8732
rect 7269 8730 7325 8732
rect 7349 8730 7405 8732
rect 7429 8730 7485 8732
rect 7189 8678 7235 8730
rect 7235 8678 7245 8730
rect 7269 8678 7299 8730
rect 7299 8678 7311 8730
rect 7311 8678 7325 8730
rect 7349 8678 7363 8730
rect 7363 8678 7375 8730
rect 7375 8678 7405 8730
rect 7429 8678 7439 8730
rect 7439 8678 7485 8730
rect 7189 8676 7245 8678
rect 7269 8676 7325 8678
rect 7349 8676 7405 8678
rect 7429 8676 7485 8678
rect 9903 8730 9959 8732
rect 9983 8730 10039 8732
rect 10063 8730 10119 8732
rect 10143 8730 10199 8732
rect 9903 8678 9949 8730
rect 9949 8678 9959 8730
rect 9983 8678 10013 8730
rect 10013 8678 10025 8730
rect 10025 8678 10039 8730
rect 10063 8678 10077 8730
rect 10077 8678 10089 8730
rect 10089 8678 10119 8730
rect 10143 8678 10153 8730
rect 10153 8678 10199 8730
rect 9903 8676 9959 8678
rect 9983 8676 10039 8678
rect 10063 8676 10119 8678
rect 10143 8676 10199 8678
rect 11260 9274 11316 9276
rect 11340 9274 11396 9276
rect 11420 9274 11476 9276
rect 11500 9274 11556 9276
rect 11260 9222 11306 9274
rect 11306 9222 11316 9274
rect 11340 9222 11370 9274
rect 11370 9222 11382 9274
rect 11382 9222 11396 9274
rect 11420 9222 11434 9274
rect 11434 9222 11446 9274
rect 11446 9222 11476 9274
rect 11500 9222 11510 9274
rect 11510 9222 11556 9274
rect 11260 9220 11316 9222
rect 11340 9220 11396 9222
rect 11420 9220 11476 9222
rect 11500 9220 11556 9222
rect 5832 8186 5888 8188
rect 5912 8186 5968 8188
rect 5992 8186 6048 8188
rect 6072 8186 6128 8188
rect 5832 8134 5878 8186
rect 5878 8134 5888 8186
rect 5912 8134 5942 8186
rect 5942 8134 5954 8186
rect 5954 8134 5968 8186
rect 5992 8134 6006 8186
rect 6006 8134 6018 8186
rect 6018 8134 6048 8186
rect 6072 8134 6082 8186
rect 6082 8134 6128 8186
rect 5832 8132 5888 8134
rect 5912 8132 5968 8134
rect 5992 8132 6048 8134
rect 6072 8132 6128 8134
rect 5832 7098 5888 7100
rect 5912 7098 5968 7100
rect 5992 7098 6048 7100
rect 6072 7098 6128 7100
rect 5832 7046 5878 7098
rect 5878 7046 5888 7098
rect 5912 7046 5942 7098
rect 5942 7046 5954 7098
rect 5954 7046 5968 7098
rect 5992 7046 6006 7098
rect 6006 7046 6018 7098
rect 6018 7046 6048 7098
rect 6072 7046 6082 7098
rect 6082 7046 6128 7098
rect 5832 7044 5888 7046
rect 5912 7044 5968 7046
rect 5992 7044 6048 7046
rect 6072 7044 6128 7046
rect 4475 6554 4531 6556
rect 4555 6554 4611 6556
rect 4635 6554 4691 6556
rect 4715 6554 4771 6556
rect 4475 6502 4521 6554
rect 4521 6502 4531 6554
rect 4555 6502 4585 6554
rect 4585 6502 4597 6554
rect 4597 6502 4611 6554
rect 4635 6502 4649 6554
rect 4649 6502 4661 6554
rect 4661 6502 4691 6554
rect 4715 6502 4725 6554
rect 4725 6502 4771 6554
rect 4475 6500 4531 6502
rect 4555 6500 4611 6502
rect 4635 6500 4691 6502
rect 4715 6500 4771 6502
rect 7189 7642 7245 7644
rect 7269 7642 7325 7644
rect 7349 7642 7405 7644
rect 7429 7642 7485 7644
rect 7189 7590 7235 7642
rect 7235 7590 7245 7642
rect 7269 7590 7299 7642
rect 7299 7590 7311 7642
rect 7311 7590 7325 7642
rect 7349 7590 7363 7642
rect 7363 7590 7375 7642
rect 7375 7590 7405 7642
rect 7429 7590 7439 7642
rect 7439 7590 7485 7642
rect 7189 7588 7245 7590
rect 7269 7588 7325 7590
rect 7349 7588 7405 7590
rect 7429 7588 7485 7590
rect 8546 8186 8602 8188
rect 8626 8186 8682 8188
rect 8706 8186 8762 8188
rect 8786 8186 8842 8188
rect 8546 8134 8592 8186
rect 8592 8134 8602 8186
rect 8626 8134 8656 8186
rect 8656 8134 8668 8186
rect 8668 8134 8682 8186
rect 8706 8134 8720 8186
rect 8720 8134 8732 8186
rect 8732 8134 8762 8186
rect 8786 8134 8796 8186
rect 8796 8134 8842 8186
rect 8546 8132 8602 8134
rect 8626 8132 8682 8134
rect 8706 8132 8762 8134
rect 8786 8132 8842 8134
rect 5832 6010 5888 6012
rect 5912 6010 5968 6012
rect 5992 6010 6048 6012
rect 6072 6010 6128 6012
rect 5832 5958 5878 6010
rect 5878 5958 5888 6010
rect 5912 5958 5942 6010
rect 5942 5958 5954 6010
rect 5954 5958 5968 6010
rect 5992 5958 6006 6010
rect 6006 5958 6018 6010
rect 6018 5958 6048 6010
rect 6072 5958 6082 6010
rect 6082 5958 6128 6010
rect 5832 5956 5888 5958
rect 5912 5956 5968 5958
rect 5992 5956 6048 5958
rect 6072 5956 6128 5958
rect 4475 5466 4531 5468
rect 4555 5466 4611 5468
rect 4635 5466 4691 5468
rect 4715 5466 4771 5468
rect 4475 5414 4521 5466
rect 4521 5414 4531 5466
rect 4555 5414 4585 5466
rect 4585 5414 4597 5466
rect 4597 5414 4611 5466
rect 4635 5414 4649 5466
rect 4649 5414 4661 5466
rect 4661 5414 4691 5466
rect 4715 5414 4725 5466
rect 4725 5414 4771 5466
rect 4475 5412 4531 5414
rect 4555 5412 4611 5414
rect 4635 5412 4691 5414
rect 4715 5412 4771 5414
rect 5832 4922 5888 4924
rect 5912 4922 5968 4924
rect 5992 4922 6048 4924
rect 6072 4922 6128 4924
rect 5832 4870 5878 4922
rect 5878 4870 5888 4922
rect 5912 4870 5942 4922
rect 5942 4870 5954 4922
rect 5954 4870 5968 4922
rect 5992 4870 6006 4922
rect 6006 4870 6018 4922
rect 6018 4870 6048 4922
rect 6072 4870 6082 4922
rect 6082 4870 6128 4922
rect 5832 4868 5888 4870
rect 5912 4868 5968 4870
rect 5992 4868 6048 4870
rect 6072 4868 6128 4870
rect 4475 4378 4531 4380
rect 4555 4378 4611 4380
rect 4635 4378 4691 4380
rect 4715 4378 4771 4380
rect 4475 4326 4521 4378
rect 4521 4326 4531 4378
rect 4555 4326 4585 4378
rect 4585 4326 4597 4378
rect 4597 4326 4611 4378
rect 4635 4326 4649 4378
rect 4649 4326 4661 4378
rect 4661 4326 4691 4378
rect 4715 4326 4725 4378
rect 4725 4326 4771 4378
rect 4475 4324 4531 4326
rect 4555 4324 4611 4326
rect 4635 4324 4691 4326
rect 4715 4324 4771 4326
rect 4475 3290 4531 3292
rect 4555 3290 4611 3292
rect 4635 3290 4691 3292
rect 4715 3290 4771 3292
rect 4475 3238 4521 3290
rect 4521 3238 4531 3290
rect 4555 3238 4585 3290
rect 4585 3238 4597 3290
rect 4597 3238 4611 3290
rect 4635 3238 4649 3290
rect 4649 3238 4661 3290
rect 4661 3238 4691 3290
rect 4715 3238 4725 3290
rect 4725 3238 4771 3290
rect 4475 3236 4531 3238
rect 4555 3236 4611 3238
rect 4635 3236 4691 3238
rect 4715 3236 4771 3238
rect 4475 2202 4531 2204
rect 4555 2202 4611 2204
rect 4635 2202 4691 2204
rect 4715 2202 4771 2204
rect 4475 2150 4521 2202
rect 4521 2150 4531 2202
rect 4555 2150 4585 2202
rect 4585 2150 4597 2202
rect 4597 2150 4611 2202
rect 4635 2150 4649 2202
rect 4649 2150 4661 2202
rect 4661 2150 4691 2202
rect 4715 2150 4725 2202
rect 4725 2150 4771 2202
rect 4475 2148 4531 2150
rect 4555 2148 4611 2150
rect 4635 2148 4691 2150
rect 4715 2148 4771 2150
rect 5832 3834 5888 3836
rect 5912 3834 5968 3836
rect 5992 3834 6048 3836
rect 6072 3834 6128 3836
rect 5832 3782 5878 3834
rect 5878 3782 5888 3834
rect 5912 3782 5942 3834
rect 5942 3782 5954 3834
rect 5954 3782 5968 3834
rect 5992 3782 6006 3834
rect 6006 3782 6018 3834
rect 6018 3782 6048 3834
rect 6072 3782 6082 3834
rect 6082 3782 6128 3834
rect 5832 3780 5888 3782
rect 5912 3780 5968 3782
rect 5992 3780 6048 3782
rect 6072 3780 6128 3782
rect 5832 2746 5888 2748
rect 5912 2746 5968 2748
rect 5992 2746 6048 2748
rect 6072 2746 6128 2748
rect 5832 2694 5878 2746
rect 5878 2694 5888 2746
rect 5912 2694 5942 2746
rect 5942 2694 5954 2746
rect 5954 2694 5968 2746
rect 5992 2694 6006 2746
rect 6006 2694 6018 2746
rect 6018 2694 6048 2746
rect 6072 2694 6082 2746
rect 6082 2694 6128 2746
rect 5832 2692 5888 2694
rect 5912 2692 5968 2694
rect 5992 2692 6048 2694
rect 6072 2692 6128 2694
rect 7189 6554 7245 6556
rect 7269 6554 7325 6556
rect 7349 6554 7405 6556
rect 7429 6554 7485 6556
rect 7189 6502 7235 6554
rect 7235 6502 7245 6554
rect 7269 6502 7299 6554
rect 7299 6502 7311 6554
rect 7311 6502 7325 6554
rect 7349 6502 7363 6554
rect 7363 6502 7375 6554
rect 7375 6502 7405 6554
rect 7429 6502 7439 6554
rect 7439 6502 7485 6554
rect 7189 6500 7245 6502
rect 7269 6500 7325 6502
rect 7349 6500 7405 6502
rect 7429 6500 7485 6502
rect 7562 6024 7618 6080
rect 7189 5466 7245 5468
rect 7269 5466 7325 5468
rect 7349 5466 7405 5468
rect 7429 5466 7485 5468
rect 7189 5414 7235 5466
rect 7235 5414 7245 5466
rect 7269 5414 7299 5466
rect 7299 5414 7311 5466
rect 7311 5414 7325 5466
rect 7349 5414 7363 5466
rect 7363 5414 7375 5466
rect 7375 5414 7405 5466
rect 7429 5414 7439 5466
rect 7439 5414 7485 5466
rect 7189 5412 7245 5414
rect 7269 5412 7325 5414
rect 7349 5412 7405 5414
rect 7429 5412 7485 5414
rect 8546 7098 8602 7100
rect 8626 7098 8682 7100
rect 8706 7098 8762 7100
rect 8786 7098 8842 7100
rect 8546 7046 8592 7098
rect 8592 7046 8602 7098
rect 8626 7046 8656 7098
rect 8656 7046 8668 7098
rect 8668 7046 8682 7098
rect 8706 7046 8720 7098
rect 8720 7046 8732 7098
rect 8732 7046 8762 7098
rect 8786 7046 8796 7098
rect 8796 7046 8842 7098
rect 8546 7044 8602 7046
rect 8626 7044 8682 7046
rect 8706 7044 8762 7046
rect 8786 7044 8842 7046
rect 11260 8186 11316 8188
rect 11340 8186 11396 8188
rect 11420 8186 11476 8188
rect 11500 8186 11556 8188
rect 11260 8134 11306 8186
rect 11306 8134 11316 8186
rect 11340 8134 11370 8186
rect 11370 8134 11382 8186
rect 11382 8134 11396 8186
rect 11420 8134 11434 8186
rect 11434 8134 11446 8186
rect 11446 8134 11476 8186
rect 11500 8134 11510 8186
rect 11510 8134 11556 8186
rect 11260 8132 11316 8134
rect 11340 8132 11396 8134
rect 11420 8132 11476 8134
rect 11500 8132 11556 8134
rect 9903 7642 9959 7644
rect 9983 7642 10039 7644
rect 10063 7642 10119 7644
rect 10143 7642 10199 7644
rect 9903 7590 9949 7642
rect 9949 7590 9959 7642
rect 9983 7590 10013 7642
rect 10013 7590 10025 7642
rect 10025 7590 10039 7642
rect 10063 7590 10077 7642
rect 10077 7590 10089 7642
rect 10089 7590 10119 7642
rect 10143 7590 10153 7642
rect 10153 7590 10199 7642
rect 9903 7588 9959 7590
rect 9983 7588 10039 7590
rect 10063 7588 10119 7590
rect 10143 7588 10199 7590
rect 11058 7384 11114 7440
rect 11260 7098 11316 7100
rect 11340 7098 11396 7100
rect 11420 7098 11476 7100
rect 11500 7098 11556 7100
rect 11260 7046 11306 7098
rect 11306 7046 11316 7098
rect 11340 7046 11370 7098
rect 11370 7046 11382 7098
rect 11382 7046 11396 7098
rect 11420 7046 11434 7098
rect 11434 7046 11446 7098
rect 11446 7046 11476 7098
rect 11500 7046 11510 7098
rect 11510 7046 11556 7098
rect 11260 7044 11316 7046
rect 11340 7044 11396 7046
rect 11420 7044 11476 7046
rect 11500 7044 11556 7046
rect 8546 6010 8602 6012
rect 8626 6010 8682 6012
rect 8706 6010 8762 6012
rect 8786 6010 8842 6012
rect 8546 5958 8592 6010
rect 8592 5958 8602 6010
rect 8626 5958 8656 6010
rect 8656 5958 8668 6010
rect 8668 5958 8682 6010
rect 8706 5958 8720 6010
rect 8720 5958 8732 6010
rect 8732 5958 8762 6010
rect 8786 5958 8796 6010
rect 8796 5958 8842 6010
rect 8546 5956 8602 5958
rect 8626 5956 8682 5958
rect 8706 5956 8762 5958
rect 8786 5956 8842 5958
rect 7189 4378 7245 4380
rect 7269 4378 7325 4380
rect 7349 4378 7405 4380
rect 7429 4378 7485 4380
rect 7189 4326 7235 4378
rect 7235 4326 7245 4378
rect 7269 4326 7299 4378
rect 7299 4326 7311 4378
rect 7311 4326 7325 4378
rect 7349 4326 7363 4378
rect 7363 4326 7375 4378
rect 7375 4326 7405 4378
rect 7429 4326 7439 4378
rect 7439 4326 7485 4378
rect 7189 4324 7245 4326
rect 7269 4324 7325 4326
rect 7349 4324 7405 4326
rect 7429 4324 7485 4326
rect 7189 3290 7245 3292
rect 7269 3290 7325 3292
rect 7349 3290 7405 3292
rect 7429 3290 7485 3292
rect 7189 3238 7235 3290
rect 7235 3238 7245 3290
rect 7269 3238 7299 3290
rect 7299 3238 7311 3290
rect 7311 3238 7325 3290
rect 7349 3238 7363 3290
rect 7363 3238 7375 3290
rect 7375 3238 7405 3290
rect 7429 3238 7439 3290
rect 7439 3238 7485 3290
rect 7189 3236 7245 3238
rect 7269 3236 7325 3238
rect 7349 3236 7405 3238
rect 7429 3236 7485 3238
rect 8546 4922 8602 4924
rect 8626 4922 8682 4924
rect 8706 4922 8762 4924
rect 8786 4922 8842 4924
rect 8546 4870 8592 4922
rect 8592 4870 8602 4922
rect 8626 4870 8656 4922
rect 8656 4870 8668 4922
rect 8668 4870 8682 4922
rect 8706 4870 8720 4922
rect 8720 4870 8732 4922
rect 8732 4870 8762 4922
rect 8786 4870 8796 4922
rect 8796 4870 8842 4922
rect 8546 4868 8602 4870
rect 8626 4868 8682 4870
rect 8706 4868 8762 4870
rect 8786 4868 8842 4870
rect 9903 6554 9959 6556
rect 9983 6554 10039 6556
rect 10063 6554 10119 6556
rect 10143 6554 10199 6556
rect 9903 6502 9949 6554
rect 9949 6502 9959 6554
rect 9983 6502 10013 6554
rect 10013 6502 10025 6554
rect 10025 6502 10039 6554
rect 10063 6502 10077 6554
rect 10077 6502 10089 6554
rect 10089 6502 10119 6554
rect 10143 6502 10153 6554
rect 10153 6502 10199 6554
rect 9903 6500 9959 6502
rect 9983 6500 10039 6502
rect 10063 6500 10119 6502
rect 10143 6500 10199 6502
rect 8546 3834 8602 3836
rect 8626 3834 8682 3836
rect 8706 3834 8762 3836
rect 8786 3834 8842 3836
rect 8546 3782 8592 3834
rect 8592 3782 8602 3834
rect 8626 3782 8656 3834
rect 8656 3782 8668 3834
rect 8668 3782 8682 3834
rect 8706 3782 8720 3834
rect 8720 3782 8732 3834
rect 8732 3782 8762 3834
rect 8786 3782 8796 3834
rect 8796 3782 8842 3834
rect 8546 3780 8602 3782
rect 8626 3780 8682 3782
rect 8706 3780 8762 3782
rect 8786 3780 8842 3782
rect 3118 1658 3174 1660
rect 3198 1658 3254 1660
rect 3278 1658 3334 1660
rect 3358 1658 3414 1660
rect 3118 1606 3164 1658
rect 3164 1606 3174 1658
rect 3198 1606 3228 1658
rect 3228 1606 3240 1658
rect 3240 1606 3254 1658
rect 3278 1606 3292 1658
rect 3292 1606 3304 1658
rect 3304 1606 3334 1658
rect 3358 1606 3368 1658
rect 3368 1606 3414 1658
rect 3118 1604 3174 1606
rect 3198 1604 3254 1606
rect 3278 1604 3334 1606
rect 3358 1604 3414 1606
rect 7189 2202 7245 2204
rect 7269 2202 7325 2204
rect 7349 2202 7405 2204
rect 7429 2202 7485 2204
rect 7189 2150 7235 2202
rect 7235 2150 7245 2202
rect 7269 2150 7299 2202
rect 7299 2150 7311 2202
rect 7311 2150 7325 2202
rect 7349 2150 7363 2202
rect 7363 2150 7375 2202
rect 7375 2150 7405 2202
rect 7429 2150 7439 2202
rect 7439 2150 7485 2202
rect 7189 2148 7245 2150
rect 7269 2148 7325 2150
rect 7349 2148 7405 2150
rect 7429 2148 7485 2150
rect 8546 2746 8602 2748
rect 8626 2746 8682 2748
rect 8706 2746 8762 2748
rect 8786 2746 8842 2748
rect 8546 2694 8592 2746
rect 8592 2694 8602 2746
rect 8626 2694 8656 2746
rect 8656 2694 8668 2746
rect 8668 2694 8682 2746
rect 8706 2694 8720 2746
rect 8720 2694 8732 2746
rect 8732 2694 8762 2746
rect 8786 2694 8796 2746
rect 8796 2694 8842 2746
rect 8546 2692 8602 2694
rect 8626 2692 8682 2694
rect 8706 2692 8762 2694
rect 8786 2692 8842 2694
rect 9903 5466 9959 5468
rect 9983 5466 10039 5468
rect 10063 5466 10119 5468
rect 10143 5466 10199 5468
rect 9903 5414 9949 5466
rect 9949 5414 9959 5466
rect 9983 5414 10013 5466
rect 10013 5414 10025 5466
rect 10025 5414 10039 5466
rect 10063 5414 10077 5466
rect 10077 5414 10089 5466
rect 10089 5414 10119 5466
rect 10143 5414 10153 5466
rect 10153 5414 10199 5466
rect 9903 5412 9959 5414
rect 9983 5412 10039 5414
rect 10063 5412 10119 5414
rect 10143 5412 10199 5414
rect 11260 6010 11316 6012
rect 11340 6010 11396 6012
rect 11420 6010 11476 6012
rect 11500 6010 11556 6012
rect 11260 5958 11306 6010
rect 11306 5958 11316 6010
rect 11340 5958 11370 6010
rect 11370 5958 11382 6010
rect 11382 5958 11396 6010
rect 11420 5958 11434 6010
rect 11434 5958 11446 6010
rect 11446 5958 11476 6010
rect 11500 5958 11510 6010
rect 11510 5958 11556 6010
rect 11260 5956 11316 5958
rect 11340 5956 11396 5958
rect 11420 5956 11476 5958
rect 11500 5956 11556 5958
rect 11260 4922 11316 4924
rect 11340 4922 11396 4924
rect 11420 4922 11476 4924
rect 11500 4922 11556 4924
rect 11260 4870 11306 4922
rect 11306 4870 11316 4922
rect 11340 4870 11370 4922
rect 11370 4870 11382 4922
rect 11382 4870 11396 4922
rect 11420 4870 11434 4922
rect 11434 4870 11446 4922
rect 11446 4870 11476 4922
rect 11500 4870 11510 4922
rect 11510 4870 11556 4922
rect 11260 4868 11316 4870
rect 11340 4868 11396 4870
rect 11420 4868 11476 4870
rect 11500 4868 11556 4870
rect 9903 4378 9959 4380
rect 9983 4378 10039 4380
rect 10063 4378 10119 4380
rect 10143 4378 10199 4380
rect 9903 4326 9949 4378
rect 9949 4326 9959 4378
rect 9983 4326 10013 4378
rect 10013 4326 10025 4378
rect 10025 4326 10039 4378
rect 10063 4326 10077 4378
rect 10077 4326 10089 4378
rect 10089 4326 10119 4378
rect 10143 4326 10153 4378
rect 10153 4326 10199 4378
rect 9903 4324 9959 4326
rect 9983 4324 10039 4326
rect 10063 4324 10119 4326
rect 10143 4324 10199 4326
rect 11260 3834 11316 3836
rect 11340 3834 11396 3836
rect 11420 3834 11476 3836
rect 11500 3834 11556 3836
rect 11260 3782 11306 3834
rect 11306 3782 11316 3834
rect 11340 3782 11370 3834
rect 11370 3782 11382 3834
rect 11382 3782 11396 3834
rect 11420 3782 11434 3834
rect 11434 3782 11446 3834
rect 11446 3782 11476 3834
rect 11500 3782 11510 3834
rect 11510 3782 11556 3834
rect 11260 3780 11316 3782
rect 11340 3780 11396 3782
rect 11420 3780 11476 3782
rect 11500 3780 11556 3782
rect 9903 3290 9959 3292
rect 9983 3290 10039 3292
rect 10063 3290 10119 3292
rect 10143 3290 10199 3292
rect 9903 3238 9949 3290
rect 9949 3238 9959 3290
rect 9983 3238 10013 3290
rect 10013 3238 10025 3290
rect 10025 3238 10039 3290
rect 10063 3238 10077 3290
rect 10077 3238 10089 3290
rect 10089 3238 10119 3290
rect 10143 3238 10153 3290
rect 10153 3238 10199 3290
rect 9903 3236 9959 3238
rect 9983 3236 10039 3238
rect 10063 3236 10119 3238
rect 10143 3236 10199 3238
rect 5832 1658 5888 1660
rect 5912 1658 5968 1660
rect 5992 1658 6048 1660
rect 6072 1658 6128 1660
rect 5832 1606 5878 1658
rect 5878 1606 5888 1658
rect 5912 1606 5942 1658
rect 5942 1606 5954 1658
rect 5954 1606 5968 1658
rect 5992 1606 6006 1658
rect 6006 1606 6018 1658
rect 6018 1606 6048 1658
rect 6072 1606 6082 1658
rect 6082 1606 6128 1658
rect 5832 1604 5888 1606
rect 5912 1604 5968 1606
rect 5992 1604 6048 1606
rect 6072 1604 6128 1606
rect 11260 2746 11316 2748
rect 11340 2746 11396 2748
rect 11420 2746 11476 2748
rect 11500 2746 11556 2748
rect 11260 2694 11306 2746
rect 11306 2694 11316 2746
rect 11340 2694 11370 2746
rect 11370 2694 11382 2746
rect 11382 2694 11396 2746
rect 11420 2694 11434 2746
rect 11434 2694 11446 2746
rect 11446 2694 11476 2746
rect 11500 2694 11510 2746
rect 11510 2694 11556 2746
rect 11260 2692 11316 2694
rect 11340 2692 11396 2694
rect 11420 2692 11476 2694
rect 11500 2692 11556 2694
rect 9903 2202 9959 2204
rect 9983 2202 10039 2204
rect 10063 2202 10119 2204
rect 10143 2202 10199 2204
rect 9903 2150 9949 2202
rect 9949 2150 9959 2202
rect 9983 2150 10013 2202
rect 10013 2150 10025 2202
rect 10025 2150 10039 2202
rect 10063 2150 10077 2202
rect 10077 2150 10089 2202
rect 10089 2150 10119 2202
rect 10143 2150 10153 2202
rect 10153 2150 10199 2202
rect 9903 2148 9959 2150
rect 9983 2148 10039 2150
rect 10063 2148 10119 2150
rect 10143 2148 10199 2150
rect 1761 1114 1817 1116
rect 1841 1114 1897 1116
rect 1921 1114 1977 1116
rect 2001 1114 2057 1116
rect 1761 1062 1807 1114
rect 1807 1062 1817 1114
rect 1841 1062 1871 1114
rect 1871 1062 1883 1114
rect 1883 1062 1897 1114
rect 1921 1062 1935 1114
rect 1935 1062 1947 1114
rect 1947 1062 1977 1114
rect 2001 1062 2011 1114
rect 2011 1062 2057 1114
rect 1761 1060 1817 1062
rect 1841 1060 1897 1062
rect 1921 1060 1977 1062
rect 2001 1060 2057 1062
rect 4475 1114 4531 1116
rect 4555 1114 4611 1116
rect 4635 1114 4691 1116
rect 4715 1114 4771 1116
rect 4475 1062 4521 1114
rect 4521 1062 4531 1114
rect 4555 1062 4585 1114
rect 4585 1062 4597 1114
rect 4597 1062 4611 1114
rect 4635 1062 4649 1114
rect 4649 1062 4661 1114
rect 4661 1062 4691 1114
rect 4715 1062 4725 1114
rect 4725 1062 4771 1114
rect 4475 1060 4531 1062
rect 4555 1060 4611 1062
rect 4635 1060 4691 1062
rect 4715 1060 4771 1062
rect 8546 1658 8602 1660
rect 8626 1658 8682 1660
rect 8706 1658 8762 1660
rect 8786 1658 8842 1660
rect 8546 1606 8592 1658
rect 8592 1606 8602 1658
rect 8626 1606 8656 1658
rect 8656 1606 8668 1658
rect 8668 1606 8682 1658
rect 8706 1606 8720 1658
rect 8720 1606 8732 1658
rect 8732 1606 8762 1658
rect 8786 1606 8796 1658
rect 8796 1606 8842 1658
rect 8546 1604 8602 1606
rect 8626 1604 8682 1606
rect 8706 1604 8762 1606
rect 8786 1604 8842 1606
rect 11260 1658 11316 1660
rect 11340 1658 11396 1660
rect 11420 1658 11476 1660
rect 11500 1658 11556 1660
rect 11260 1606 11306 1658
rect 11306 1606 11316 1658
rect 11340 1606 11370 1658
rect 11370 1606 11382 1658
rect 11382 1606 11396 1658
rect 11420 1606 11434 1658
rect 11434 1606 11446 1658
rect 11446 1606 11476 1658
rect 11500 1606 11510 1658
rect 11510 1606 11556 1658
rect 11260 1604 11316 1606
rect 11340 1604 11396 1606
rect 11420 1604 11476 1606
rect 11500 1604 11556 1606
rect 7189 1114 7245 1116
rect 7269 1114 7325 1116
rect 7349 1114 7405 1116
rect 7429 1114 7485 1116
rect 7189 1062 7235 1114
rect 7235 1062 7245 1114
rect 7269 1062 7299 1114
rect 7299 1062 7311 1114
rect 7311 1062 7325 1114
rect 7349 1062 7363 1114
rect 7363 1062 7375 1114
rect 7375 1062 7405 1114
rect 7429 1062 7439 1114
rect 7439 1062 7485 1114
rect 7189 1060 7245 1062
rect 7269 1060 7325 1062
rect 7349 1060 7405 1062
rect 7429 1060 7485 1062
rect 9903 1114 9959 1116
rect 9983 1114 10039 1116
rect 10063 1114 10119 1116
rect 10143 1114 10199 1116
rect 9903 1062 9949 1114
rect 9949 1062 9959 1114
rect 9983 1062 10013 1114
rect 10013 1062 10025 1114
rect 10025 1062 10039 1114
rect 10063 1062 10077 1114
rect 10077 1062 10089 1114
rect 10089 1062 10119 1114
rect 10143 1062 10153 1114
rect 10153 1062 10199 1114
rect 9903 1060 9959 1062
rect 9983 1060 10039 1062
rect 10063 1060 10119 1062
rect 10143 1060 10199 1062
rect 3118 570 3174 572
rect 3198 570 3254 572
rect 3278 570 3334 572
rect 3358 570 3414 572
rect 3118 518 3164 570
rect 3164 518 3174 570
rect 3198 518 3228 570
rect 3228 518 3240 570
rect 3240 518 3254 570
rect 3278 518 3292 570
rect 3292 518 3304 570
rect 3304 518 3334 570
rect 3358 518 3368 570
rect 3368 518 3414 570
rect 3118 516 3174 518
rect 3198 516 3254 518
rect 3278 516 3334 518
rect 3358 516 3414 518
rect 5832 570 5888 572
rect 5912 570 5968 572
rect 5992 570 6048 572
rect 6072 570 6128 572
rect 5832 518 5878 570
rect 5878 518 5888 570
rect 5912 518 5942 570
rect 5942 518 5954 570
rect 5954 518 5968 570
rect 5992 518 6006 570
rect 6006 518 6018 570
rect 6018 518 6048 570
rect 6072 518 6082 570
rect 6082 518 6128 570
rect 5832 516 5888 518
rect 5912 516 5968 518
rect 5992 516 6048 518
rect 6072 516 6128 518
rect 8546 570 8602 572
rect 8626 570 8682 572
rect 8706 570 8762 572
rect 8786 570 8842 572
rect 8546 518 8592 570
rect 8592 518 8602 570
rect 8626 518 8656 570
rect 8656 518 8668 570
rect 8668 518 8682 570
rect 8706 518 8720 570
rect 8720 518 8732 570
rect 8732 518 8762 570
rect 8786 518 8796 570
rect 8796 518 8842 570
rect 8546 516 8602 518
rect 8626 516 8682 518
rect 8706 516 8762 518
rect 8786 516 8842 518
rect 11260 570 11316 572
rect 11340 570 11396 572
rect 11420 570 11476 572
rect 11500 570 11556 572
rect 11260 518 11306 570
rect 11306 518 11316 570
rect 11340 518 11370 570
rect 11370 518 11382 570
rect 11382 518 11396 570
rect 11420 518 11434 570
rect 11434 518 11446 570
rect 11446 518 11476 570
rect 11500 518 11510 570
rect 11510 518 11556 570
rect 11260 516 11316 518
rect 11340 516 11396 518
rect 11420 516 11476 518
rect 11500 516 11556 518
<< metal3 >>
rect 3108 9280 3424 9281
rect 3108 9216 3114 9280
rect 3178 9216 3194 9280
rect 3258 9216 3274 9280
rect 3338 9216 3354 9280
rect 3418 9216 3424 9280
rect 3108 9215 3424 9216
rect 5822 9280 6138 9281
rect 5822 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5988 9280
rect 6052 9216 6068 9280
rect 6132 9216 6138 9280
rect 5822 9215 6138 9216
rect 8536 9280 8852 9281
rect 8536 9216 8542 9280
rect 8606 9216 8622 9280
rect 8686 9216 8702 9280
rect 8766 9216 8782 9280
rect 8846 9216 8852 9280
rect 8536 9215 8852 9216
rect 11250 9280 11566 9281
rect 11250 9216 11256 9280
rect 11320 9216 11336 9280
rect 11400 9216 11416 9280
rect 11480 9216 11496 9280
rect 11560 9216 11566 9280
rect 11250 9215 11566 9216
rect 1751 8736 2067 8737
rect 1751 8672 1757 8736
rect 1821 8672 1837 8736
rect 1901 8672 1917 8736
rect 1981 8672 1997 8736
rect 2061 8672 2067 8736
rect 1751 8671 2067 8672
rect 4465 8736 4781 8737
rect 4465 8672 4471 8736
rect 4535 8672 4551 8736
rect 4615 8672 4631 8736
rect 4695 8672 4711 8736
rect 4775 8672 4781 8736
rect 4465 8671 4781 8672
rect 7179 8736 7495 8737
rect 7179 8672 7185 8736
rect 7249 8672 7265 8736
rect 7329 8672 7345 8736
rect 7409 8672 7425 8736
rect 7489 8672 7495 8736
rect 7179 8671 7495 8672
rect 9893 8736 10209 8737
rect 9893 8672 9899 8736
rect 9963 8672 9979 8736
rect 10043 8672 10059 8736
rect 10123 8672 10139 8736
rect 10203 8672 10209 8736
rect 9893 8671 10209 8672
rect 3108 8192 3424 8193
rect 3108 8128 3114 8192
rect 3178 8128 3194 8192
rect 3258 8128 3274 8192
rect 3338 8128 3354 8192
rect 3418 8128 3424 8192
rect 3108 8127 3424 8128
rect 5822 8192 6138 8193
rect 5822 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5988 8192
rect 6052 8128 6068 8192
rect 6132 8128 6138 8192
rect 5822 8127 6138 8128
rect 8536 8192 8852 8193
rect 8536 8128 8542 8192
rect 8606 8128 8622 8192
rect 8686 8128 8702 8192
rect 8766 8128 8782 8192
rect 8846 8128 8852 8192
rect 8536 8127 8852 8128
rect 11250 8192 11566 8193
rect 11250 8128 11256 8192
rect 11320 8128 11336 8192
rect 11400 8128 11416 8192
rect 11480 8128 11496 8192
rect 11560 8128 11566 8192
rect 11250 8127 11566 8128
rect 1751 7648 2067 7649
rect 1751 7584 1757 7648
rect 1821 7584 1837 7648
rect 1901 7584 1917 7648
rect 1981 7584 1997 7648
rect 2061 7584 2067 7648
rect 1751 7583 2067 7584
rect 4465 7648 4781 7649
rect 4465 7584 4471 7648
rect 4535 7584 4551 7648
rect 4615 7584 4631 7648
rect 4695 7584 4711 7648
rect 4775 7584 4781 7648
rect 4465 7583 4781 7584
rect 7179 7648 7495 7649
rect 7179 7584 7185 7648
rect 7249 7584 7265 7648
rect 7329 7584 7345 7648
rect 7409 7584 7425 7648
rect 7489 7584 7495 7648
rect 7179 7583 7495 7584
rect 9893 7648 10209 7649
rect 9893 7584 9899 7648
rect 9963 7584 9979 7648
rect 10043 7584 10059 7648
rect 10123 7584 10139 7648
rect 10203 7584 10209 7648
rect 9893 7583 10209 7584
rect 11053 7442 11119 7445
rect 11600 7442 12000 7472
rect 11053 7440 12000 7442
rect 11053 7384 11058 7440
rect 11114 7384 12000 7440
rect 11053 7382 12000 7384
rect 11053 7379 11119 7382
rect 11600 7352 12000 7382
rect 3108 7104 3424 7105
rect 3108 7040 3114 7104
rect 3178 7040 3194 7104
rect 3258 7040 3274 7104
rect 3338 7040 3354 7104
rect 3418 7040 3424 7104
rect 3108 7039 3424 7040
rect 5822 7104 6138 7105
rect 5822 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5988 7104
rect 6052 7040 6068 7104
rect 6132 7040 6138 7104
rect 5822 7039 6138 7040
rect 8536 7104 8852 7105
rect 8536 7040 8542 7104
rect 8606 7040 8622 7104
rect 8686 7040 8702 7104
rect 8766 7040 8782 7104
rect 8846 7040 8852 7104
rect 8536 7039 8852 7040
rect 11250 7104 11566 7105
rect 11250 7040 11256 7104
rect 11320 7040 11336 7104
rect 11400 7040 11416 7104
rect 11480 7040 11496 7104
rect 11560 7040 11566 7104
rect 11250 7039 11566 7040
rect 1751 6560 2067 6561
rect 1751 6496 1757 6560
rect 1821 6496 1837 6560
rect 1901 6496 1917 6560
rect 1981 6496 1997 6560
rect 2061 6496 2067 6560
rect 1751 6495 2067 6496
rect 4465 6560 4781 6561
rect 4465 6496 4471 6560
rect 4535 6496 4551 6560
rect 4615 6496 4631 6560
rect 4695 6496 4711 6560
rect 4775 6496 4781 6560
rect 4465 6495 4781 6496
rect 7179 6560 7495 6561
rect 7179 6496 7185 6560
rect 7249 6496 7265 6560
rect 7329 6496 7345 6560
rect 7409 6496 7425 6560
rect 7489 6496 7495 6560
rect 7179 6495 7495 6496
rect 9893 6560 10209 6561
rect 9893 6496 9899 6560
rect 9963 6496 9979 6560
rect 10043 6496 10059 6560
rect 10123 6496 10139 6560
rect 10203 6496 10209 6560
rect 9893 6495 10209 6496
rect 7557 6084 7623 6085
rect 7557 6082 7604 6084
rect 7512 6080 7604 6082
rect 7512 6024 7562 6080
rect 7512 6022 7604 6024
rect 7557 6020 7604 6022
rect 7668 6020 7674 6084
rect 7557 6019 7623 6020
rect 3108 6016 3424 6017
rect 3108 5952 3114 6016
rect 3178 5952 3194 6016
rect 3258 5952 3274 6016
rect 3338 5952 3354 6016
rect 3418 5952 3424 6016
rect 3108 5951 3424 5952
rect 5822 6016 6138 6017
rect 5822 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5988 6016
rect 6052 5952 6068 6016
rect 6132 5952 6138 6016
rect 5822 5951 6138 5952
rect 8536 6016 8852 6017
rect 8536 5952 8542 6016
rect 8606 5952 8622 6016
rect 8686 5952 8702 6016
rect 8766 5952 8782 6016
rect 8846 5952 8852 6016
rect 8536 5951 8852 5952
rect 11250 6016 11566 6017
rect 11250 5952 11256 6016
rect 11320 5952 11336 6016
rect 11400 5952 11416 6016
rect 11480 5952 11496 6016
rect 11560 5952 11566 6016
rect 11250 5951 11566 5952
rect 1751 5472 2067 5473
rect 1751 5408 1757 5472
rect 1821 5408 1837 5472
rect 1901 5408 1917 5472
rect 1981 5408 1997 5472
rect 2061 5408 2067 5472
rect 1751 5407 2067 5408
rect 4465 5472 4781 5473
rect 4465 5408 4471 5472
rect 4535 5408 4551 5472
rect 4615 5408 4631 5472
rect 4695 5408 4711 5472
rect 4775 5408 4781 5472
rect 4465 5407 4781 5408
rect 7179 5472 7495 5473
rect 7179 5408 7185 5472
rect 7249 5408 7265 5472
rect 7329 5408 7345 5472
rect 7409 5408 7425 5472
rect 7489 5408 7495 5472
rect 7179 5407 7495 5408
rect 9893 5472 10209 5473
rect 9893 5408 9899 5472
rect 9963 5408 9979 5472
rect 10043 5408 10059 5472
rect 10123 5408 10139 5472
rect 10203 5408 10209 5472
rect 9893 5407 10209 5408
rect 3108 4928 3424 4929
rect 3108 4864 3114 4928
rect 3178 4864 3194 4928
rect 3258 4864 3274 4928
rect 3338 4864 3354 4928
rect 3418 4864 3424 4928
rect 3108 4863 3424 4864
rect 5822 4928 6138 4929
rect 5822 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5988 4928
rect 6052 4864 6068 4928
rect 6132 4864 6138 4928
rect 5822 4863 6138 4864
rect 8536 4928 8852 4929
rect 8536 4864 8542 4928
rect 8606 4864 8622 4928
rect 8686 4864 8702 4928
rect 8766 4864 8782 4928
rect 8846 4864 8852 4928
rect 8536 4863 8852 4864
rect 11250 4928 11566 4929
rect 11250 4864 11256 4928
rect 11320 4864 11336 4928
rect 11400 4864 11416 4928
rect 11480 4864 11496 4928
rect 11560 4864 11566 4928
rect 11250 4863 11566 4864
rect 1751 4384 2067 4385
rect 1751 4320 1757 4384
rect 1821 4320 1837 4384
rect 1901 4320 1917 4384
rect 1981 4320 1997 4384
rect 2061 4320 2067 4384
rect 1751 4319 2067 4320
rect 4465 4384 4781 4385
rect 4465 4320 4471 4384
rect 4535 4320 4551 4384
rect 4615 4320 4631 4384
rect 4695 4320 4711 4384
rect 4775 4320 4781 4384
rect 4465 4319 4781 4320
rect 7179 4384 7495 4385
rect 7179 4320 7185 4384
rect 7249 4320 7265 4384
rect 7329 4320 7345 4384
rect 7409 4320 7425 4384
rect 7489 4320 7495 4384
rect 7179 4319 7495 4320
rect 9893 4384 10209 4385
rect 9893 4320 9899 4384
rect 9963 4320 9979 4384
rect 10043 4320 10059 4384
rect 10123 4320 10139 4384
rect 10203 4320 10209 4384
rect 9893 4319 10209 4320
rect 3108 3840 3424 3841
rect 3108 3776 3114 3840
rect 3178 3776 3194 3840
rect 3258 3776 3274 3840
rect 3338 3776 3354 3840
rect 3418 3776 3424 3840
rect 3108 3775 3424 3776
rect 5822 3840 6138 3841
rect 5822 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5988 3840
rect 6052 3776 6068 3840
rect 6132 3776 6138 3840
rect 5822 3775 6138 3776
rect 8536 3840 8852 3841
rect 8536 3776 8542 3840
rect 8606 3776 8622 3840
rect 8686 3776 8702 3840
rect 8766 3776 8782 3840
rect 8846 3776 8852 3840
rect 8536 3775 8852 3776
rect 11250 3840 11566 3841
rect 11250 3776 11256 3840
rect 11320 3776 11336 3840
rect 11400 3776 11416 3840
rect 11480 3776 11496 3840
rect 11560 3776 11566 3840
rect 11250 3775 11566 3776
rect 1751 3296 2067 3297
rect 1751 3232 1757 3296
rect 1821 3232 1837 3296
rect 1901 3232 1917 3296
rect 1981 3232 1997 3296
rect 2061 3232 2067 3296
rect 1751 3231 2067 3232
rect 4465 3296 4781 3297
rect 4465 3232 4471 3296
rect 4535 3232 4551 3296
rect 4615 3232 4631 3296
rect 4695 3232 4711 3296
rect 4775 3232 4781 3296
rect 4465 3231 4781 3232
rect 7179 3296 7495 3297
rect 7179 3232 7185 3296
rect 7249 3232 7265 3296
rect 7329 3232 7345 3296
rect 7409 3232 7425 3296
rect 7489 3232 7495 3296
rect 7179 3231 7495 3232
rect 9893 3296 10209 3297
rect 9893 3232 9899 3296
rect 9963 3232 9979 3296
rect 10043 3232 10059 3296
rect 10123 3232 10139 3296
rect 10203 3232 10209 3296
rect 9893 3231 10209 3232
rect 3108 2752 3424 2753
rect 3108 2688 3114 2752
rect 3178 2688 3194 2752
rect 3258 2688 3274 2752
rect 3338 2688 3354 2752
rect 3418 2688 3424 2752
rect 3108 2687 3424 2688
rect 5822 2752 6138 2753
rect 5822 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5988 2752
rect 6052 2688 6068 2752
rect 6132 2688 6138 2752
rect 5822 2687 6138 2688
rect 8536 2752 8852 2753
rect 8536 2688 8542 2752
rect 8606 2688 8622 2752
rect 8686 2688 8702 2752
rect 8766 2688 8782 2752
rect 8846 2688 8852 2752
rect 8536 2687 8852 2688
rect 11250 2752 11566 2753
rect 11250 2688 11256 2752
rect 11320 2688 11336 2752
rect 11400 2688 11416 2752
rect 11480 2688 11496 2752
rect 11560 2688 11566 2752
rect 11250 2687 11566 2688
rect 7598 2484 7604 2548
rect 7668 2546 7674 2548
rect 11600 2546 12000 2576
rect 7668 2486 12000 2546
rect 7668 2484 7674 2486
rect 11600 2456 12000 2486
rect 1751 2208 2067 2209
rect 1751 2144 1757 2208
rect 1821 2144 1837 2208
rect 1901 2144 1917 2208
rect 1981 2144 1997 2208
rect 2061 2144 2067 2208
rect 1751 2143 2067 2144
rect 4465 2208 4781 2209
rect 4465 2144 4471 2208
rect 4535 2144 4551 2208
rect 4615 2144 4631 2208
rect 4695 2144 4711 2208
rect 4775 2144 4781 2208
rect 4465 2143 4781 2144
rect 7179 2208 7495 2209
rect 7179 2144 7185 2208
rect 7249 2144 7265 2208
rect 7329 2144 7345 2208
rect 7409 2144 7425 2208
rect 7489 2144 7495 2208
rect 7179 2143 7495 2144
rect 9893 2208 10209 2209
rect 9893 2144 9899 2208
rect 9963 2144 9979 2208
rect 10043 2144 10059 2208
rect 10123 2144 10139 2208
rect 10203 2144 10209 2208
rect 9893 2143 10209 2144
rect 3108 1664 3424 1665
rect 3108 1600 3114 1664
rect 3178 1600 3194 1664
rect 3258 1600 3274 1664
rect 3338 1600 3354 1664
rect 3418 1600 3424 1664
rect 3108 1599 3424 1600
rect 5822 1664 6138 1665
rect 5822 1600 5828 1664
rect 5892 1600 5908 1664
rect 5972 1600 5988 1664
rect 6052 1600 6068 1664
rect 6132 1600 6138 1664
rect 5822 1599 6138 1600
rect 8536 1664 8852 1665
rect 8536 1600 8542 1664
rect 8606 1600 8622 1664
rect 8686 1600 8702 1664
rect 8766 1600 8782 1664
rect 8846 1600 8852 1664
rect 8536 1599 8852 1600
rect 11250 1664 11566 1665
rect 11250 1600 11256 1664
rect 11320 1600 11336 1664
rect 11400 1600 11416 1664
rect 11480 1600 11496 1664
rect 11560 1600 11566 1664
rect 11250 1599 11566 1600
rect 1751 1120 2067 1121
rect 1751 1056 1757 1120
rect 1821 1056 1837 1120
rect 1901 1056 1917 1120
rect 1981 1056 1997 1120
rect 2061 1056 2067 1120
rect 1751 1055 2067 1056
rect 4465 1120 4781 1121
rect 4465 1056 4471 1120
rect 4535 1056 4551 1120
rect 4615 1056 4631 1120
rect 4695 1056 4711 1120
rect 4775 1056 4781 1120
rect 4465 1055 4781 1056
rect 7179 1120 7495 1121
rect 7179 1056 7185 1120
rect 7249 1056 7265 1120
rect 7329 1056 7345 1120
rect 7409 1056 7425 1120
rect 7489 1056 7495 1120
rect 7179 1055 7495 1056
rect 9893 1120 10209 1121
rect 9893 1056 9899 1120
rect 9963 1056 9979 1120
rect 10043 1056 10059 1120
rect 10123 1056 10139 1120
rect 10203 1056 10209 1120
rect 9893 1055 10209 1056
rect 3108 576 3424 577
rect 3108 512 3114 576
rect 3178 512 3194 576
rect 3258 512 3274 576
rect 3338 512 3354 576
rect 3418 512 3424 576
rect 3108 511 3424 512
rect 5822 576 6138 577
rect 5822 512 5828 576
rect 5892 512 5908 576
rect 5972 512 5988 576
rect 6052 512 6068 576
rect 6132 512 6138 576
rect 5822 511 6138 512
rect 8536 576 8852 577
rect 8536 512 8542 576
rect 8606 512 8622 576
rect 8686 512 8702 576
rect 8766 512 8782 576
rect 8846 512 8852 576
rect 8536 511 8852 512
rect 11250 576 11566 577
rect 11250 512 11256 576
rect 11320 512 11336 576
rect 11400 512 11416 576
rect 11480 512 11496 576
rect 11560 512 11566 576
rect 11250 511 11566 512
<< via3 >>
rect 3114 9276 3178 9280
rect 3114 9220 3118 9276
rect 3118 9220 3174 9276
rect 3174 9220 3178 9276
rect 3114 9216 3178 9220
rect 3194 9276 3258 9280
rect 3194 9220 3198 9276
rect 3198 9220 3254 9276
rect 3254 9220 3258 9276
rect 3194 9216 3258 9220
rect 3274 9276 3338 9280
rect 3274 9220 3278 9276
rect 3278 9220 3334 9276
rect 3334 9220 3338 9276
rect 3274 9216 3338 9220
rect 3354 9276 3418 9280
rect 3354 9220 3358 9276
rect 3358 9220 3414 9276
rect 3414 9220 3418 9276
rect 3354 9216 3418 9220
rect 5828 9276 5892 9280
rect 5828 9220 5832 9276
rect 5832 9220 5888 9276
rect 5888 9220 5892 9276
rect 5828 9216 5892 9220
rect 5908 9276 5972 9280
rect 5908 9220 5912 9276
rect 5912 9220 5968 9276
rect 5968 9220 5972 9276
rect 5908 9216 5972 9220
rect 5988 9276 6052 9280
rect 5988 9220 5992 9276
rect 5992 9220 6048 9276
rect 6048 9220 6052 9276
rect 5988 9216 6052 9220
rect 6068 9276 6132 9280
rect 6068 9220 6072 9276
rect 6072 9220 6128 9276
rect 6128 9220 6132 9276
rect 6068 9216 6132 9220
rect 8542 9276 8606 9280
rect 8542 9220 8546 9276
rect 8546 9220 8602 9276
rect 8602 9220 8606 9276
rect 8542 9216 8606 9220
rect 8622 9276 8686 9280
rect 8622 9220 8626 9276
rect 8626 9220 8682 9276
rect 8682 9220 8686 9276
rect 8622 9216 8686 9220
rect 8702 9276 8766 9280
rect 8702 9220 8706 9276
rect 8706 9220 8762 9276
rect 8762 9220 8766 9276
rect 8702 9216 8766 9220
rect 8782 9276 8846 9280
rect 8782 9220 8786 9276
rect 8786 9220 8842 9276
rect 8842 9220 8846 9276
rect 8782 9216 8846 9220
rect 11256 9276 11320 9280
rect 11256 9220 11260 9276
rect 11260 9220 11316 9276
rect 11316 9220 11320 9276
rect 11256 9216 11320 9220
rect 11336 9276 11400 9280
rect 11336 9220 11340 9276
rect 11340 9220 11396 9276
rect 11396 9220 11400 9276
rect 11336 9216 11400 9220
rect 11416 9276 11480 9280
rect 11416 9220 11420 9276
rect 11420 9220 11476 9276
rect 11476 9220 11480 9276
rect 11416 9216 11480 9220
rect 11496 9276 11560 9280
rect 11496 9220 11500 9276
rect 11500 9220 11556 9276
rect 11556 9220 11560 9276
rect 11496 9216 11560 9220
rect 1757 8732 1821 8736
rect 1757 8676 1761 8732
rect 1761 8676 1817 8732
rect 1817 8676 1821 8732
rect 1757 8672 1821 8676
rect 1837 8732 1901 8736
rect 1837 8676 1841 8732
rect 1841 8676 1897 8732
rect 1897 8676 1901 8732
rect 1837 8672 1901 8676
rect 1917 8732 1981 8736
rect 1917 8676 1921 8732
rect 1921 8676 1977 8732
rect 1977 8676 1981 8732
rect 1917 8672 1981 8676
rect 1997 8732 2061 8736
rect 1997 8676 2001 8732
rect 2001 8676 2057 8732
rect 2057 8676 2061 8732
rect 1997 8672 2061 8676
rect 4471 8732 4535 8736
rect 4471 8676 4475 8732
rect 4475 8676 4531 8732
rect 4531 8676 4535 8732
rect 4471 8672 4535 8676
rect 4551 8732 4615 8736
rect 4551 8676 4555 8732
rect 4555 8676 4611 8732
rect 4611 8676 4615 8732
rect 4551 8672 4615 8676
rect 4631 8732 4695 8736
rect 4631 8676 4635 8732
rect 4635 8676 4691 8732
rect 4691 8676 4695 8732
rect 4631 8672 4695 8676
rect 4711 8732 4775 8736
rect 4711 8676 4715 8732
rect 4715 8676 4771 8732
rect 4771 8676 4775 8732
rect 4711 8672 4775 8676
rect 7185 8732 7249 8736
rect 7185 8676 7189 8732
rect 7189 8676 7245 8732
rect 7245 8676 7249 8732
rect 7185 8672 7249 8676
rect 7265 8732 7329 8736
rect 7265 8676 7269 8732
rect 7269 8676 7325 8732
rect 7325 8676 7329 8732
rect 7265 8672 7329 8676
rect 7345 8732 7409 8736
rect 7345 8676 7349 8732
rect 7349 8676 7405 8732
rect 7405 8676 7409 8732
rect 7345 8672 7409 8676
rect 7425 8732 7489 8736
rect 7425 8676 7429 8732
rect 7429 8676 7485 8732
rect 7485 8676 7489 8732
rect 7425 8672 7489 8676
rect 9899 8732 9963 8736
rect 9899 8676 9903 8732
rect 9903 8676 9959 8732
rect 9959 8676 9963 8732
rect 9899 8672 9963 8676
rect 9979 8732 10043 8736
rect 9979 8676 9983 8732
rect 9983 8676 10039 8732
rect 10039 8676 10043 8732
rect 9979 8672 10043 8676
rect 10059 8732 10123 8736
rect 10059 8676 10063 8732
rect 10063 8676 10119 8732
rect 10119 8676 10123 8732
rect 10059 8672 10123 8676
rect 10139 8732 10203 8736
rect 10139 8676 10143 8732
rect 10143 8676 10199 8732
rect 10199 8676 10203 8732
rect 10139 8672 10203 8676
rect 3114 8188 3178 8192
rect 3114 8132 3118 8188
rect 3118 8132 3174 8188
rect 3174 8132 3178 8188
rect 3114 8128 3178 8132
rect 3194 8188 3258 8192
rect 3194 8132 3198 8188
rect 3198 8132 3254 8188
rect 3254 8132 3258 8188
rect 3194 8128 3258 8132
rect 3274 8188 3338 8192
rect 3274 8132 3278 8188
rect 3278 8132 3334 8188
rect 3334 8132 3338 8188
rect 3274 8128 3338 8132
rect 3354 8188 3418 8192
rect 3354 8132 3358 8188
rect 3358 8132 3414 8188
rect 3414 8132 3418 8188
rect 3354 8128 3418 8132
rect 5828 8188 5892 8192
rect 5828 8132 5832 8188
rect 5832 8132 5888 8188
rect 5888 8132 5892 8188
rect 5828 8128 5892 8132
rect 5908 8188 5972 8192
rect 5908 8132 5912 8188
rect 5912 8132 5968 8188
rect 5968 8132 5972 8188
rect 5908 8128 5972 8132
rect 5988 8188 6052 8192
rect 5988 8132 5992 8188
rect 5992 8132 6048 8188
rect 6048 8132 6052 8188
rect 5988 8128 6052 8132
rect 6068 8188 6132 8192
rect 6068 8132 6072 8188
rect 6072 8132 6128 8188
rect 6128 8132 6132 8188
rect 6068 8128 6132 8132
rect 8542 8188 8606 8192
rect 8542 8132 8546 8188
rect 8546 8132 8602 8188
rect 8602 8132 8606 8188
rect 8542 8128 8606 8132
rect 8622 8188 8686 8192
rect 8622 8132 8626 8188
rect 8626 8132 8682 8188
rect 8682 8132 8686 8188
rect 8622 8128 8686 8132
rect 8702 8188 8766 8192
rect 8702 8132 8706 8188
rect 8706 8132 8762 8188
rect 8762 8132 8766 8188
rect 8702 8128 8766 8132
rect 8782 8188 8846 8192
rect 8782 8132 8786 8188
rect 8786 8132 8842 8188
rect 8842 8132 8846 8188
rect 8782 8128 8846 8132
rect 11256 8188 11320 8192
rect 11256 8132 11260 8188
rect 11260 8132 11316 8188
rect 11316 8132 11320 8188
rect 11256 8128 11320 8132
rect 11336 8188 11400 8192
rect 11336 8132 11340 8188
rect 11340 8132 11396 8188
rect 11396 8132 11400 8188
rect 11336 8128 11400 8132
rect 11416 8188 11480 8192
rect 11416 8132 11420 8188
rect 11420 8132 11476 8188
rect 11476 8132 11480 8188
rect 11416 8128 11480 8132
rect 11496 8188 11560 8192
rect 11496 8132 11500 8188
rect 11500 8132 11556 8188
rect 11556 8132 11560 8188
rect 11496 8128 11560 8132
rect 1757 7644 1821 7648
rect 1757 7588 1761 7644
rect 1761 7588 1817 7644
rect 1817 7588 1821 7644
rect 1757 7584 1821 7588
rect 1837 7644 1901 7648
rect 1837 7588 1841 7644
rect 1841 7588 1897 7644
rect 1897 7588 1901 7644
rect 1837 7584 1901 7588
rect 1917 7644 1981 7648
rect 1917 7588 1921 7644
rect 1921 7588 1977 7644
rect 1977 7588 1981 7644
rect 1917 7584 1981 7588
rect 1997 7644 2061 7648
rect 1997 7588 2001 7644
rect 2001 7588 2057 7644
rect 2057 7588 2061 7644
rect 1997 7584 2061 7588
rect 4471 7644 4535 7648
rect 4471 7588 4475 7644
rect 4475 7588 4531 7644
rect 4531 7588 4535 7644
rect 4471 7584 4535 7588
rect 4551 7644 4615 7648
rect 4551 7588 4555 7644
rect 4555 7588 4611 7644
rect 4611 7588 4615 7644
rect 4551 7584 4615 7588
rect 4631 7644 4695 7648
rect 4631 7588 4635 7644
rect 4635 7588 4691 7644
rect 4691 7588 4695 7644
rect 4631 7584 4695 7588
rect 4711 7644 4775 7648
rect 4711 7588 4715 7644
rect 4715 7588 4771 7644
rect 4771 7588 4775 7644
rect 4711 7584 4775 7588
rect 7185 7644 7249 7648
rect 7185 7588 7189 7644
rect 7189 7588 7245 7644
rect 7245 7588 7249 7644
rect 7185 7584 7249 7588
rect 7265 7644 7329 7648
rect 7265 7588 7269 7644
rect 7269 7588 7325 7644
rect 7325 7588 7329 7644
rect 7265 7584 7329 7588
rect 7345 7644 7409 7648
rect 7345 7588 7349 7644
rect 7349 7588 7405 7644
rect 7405 7588 7409 7644
rect 7345 7584 7409 7588
rect 7425 7644 7489 7648
rect 7425 7588 7429 7644
rect 7429 7588 7485 7644
rect 7485 7588 7489 7644
rect 7425 7584 7489 7588
rect 9899 7644 9963 7648
rect 9899 7588 9903 7644
rect 9903 7588 9959 7644
rect 9959 7588 9963 7644
rect 9899 7584 9963 7588
rect 9979 7644 10043 7648
rect 9979 7588 9983 7644
rect 9983 7588 10039 7644
rect 10039 7588 10043 7644
rect 9979 7584 10043 7588
rect 10059 7644 10123 7648
rect 10059 7588 10063 7644
rect 10063 7588 10119 7644
rect 10119 7588 10123 7644
rect 10059 7584 10123 7588
rect 10139 7644 10203 7648
rect 10139 7588 10143 7644
rect 10143 7588 10199 7644
rect 10199 7588 10203 7644
rect 10139 7584 10203 7588
rect 3114 7100 3178 7104
rect 3114 7044 3118 7100
rect 3118 7044 3174 7100
rect 3174 7044 3178 7100
rect 3114 7040 3178 7044
rect 3194 7100 3258 7104
rect 3194 7044 3198 7100
rect 3198 7044 3254 7100
rect 3254 7044 3258 7100
rect 3194 7040 3258 7044
rect 3274 7100 3338 7104
rect 3274 7044 3278 7100
rect 3278 7044 3334 7100
rect 3334 7044 3338 7100
rect 3274 7040 3338 7044
rect 3354 7100 3418 7104
rect 3354 7044 3358 7100
rect 3358 7044 3414 7100
rect 3414 7044 3418 7100
rect 3354 7040 3418 7044
rect 5828 7100 5892 7104
rect 5828 7044 5832 7100
rect 5832 7044 5888 7100
rect 5888 7044 5892 7100
rect 5828 7040 5892 7044
rect 5908 7100 5972 7104
rect 5908 7044 5912 7100
rect 5912 7044 5968 7100
rect 5968 7044 5972 7100
rect 5908 7040 5972 7044
rect 5988 7100 6052 7104
rect 5988 7044 5992 7100
rect 5992 7044 6048 7100
rect 6048 7044 6052 7100
rect 5988 7040 6052 7044
rect 6068 7100 6132 7104
rect 6068 7044 6072 7100
rect 6072 7044 6128 7100
rect 6128 7044 6132 7100
rect 6068 7040 6132 7044
rect 8542 7100 8606 7104
rect 8542 7044 8546 7100
rect 8546 7044 8602 7100
rect 8602 7044 8606 7100
rect 8542 7040 8606 7044
rect 8622 7100 8686 7104
rect 8622 7044 8626 7100
rect 8626 7044 8682 7100
rect 8682 7044 8686 7100
rect 8622 7040 8686 7044
rect 8702 7100 8766 7104
rect 8702 7044 8706 7100
rect 8706 7044 8762 7100
rect 8762 7044 8766 7100
rect 8702 7040 8766 7044
rect 8782 7100 8846 7104
rect 8782 7044 8786 7100
rect 8786 7044 8842 7100
rect 8842 7044 8846 7100
rect 8782 7040 8846 7044
rect 11256 7100 11320 7104
rect 11256 7044 11260 7100
rect 11260 7044 11316 7100
rect 11316 7044 11320 7100
rect 11256 7040 11320 7044
rect 11336 7100 11400 7104
rect 11336 7044 11340 7100
rect 11340 7044 11396 7100
rect 11396 7044 11400 7100
rect 11336 7040 11400 7044
rect 11416 7100 11480 7104
rect 11416 7044 11420 7100
rect 11420 7044 11476 7100
rect 11476 7044 11480 7100
rect 11416 7040 11480 7044
rect 11496 7100 11560 7104
rect 11496 7044 11500 7100
rect 11500 7044 11556 7100
rect 11556 7044 11560 7100
rect 11496 7040 11560 7044
rect 1757 6556 1821 6560
rect 1757 6500 1761 6556
rect 1761 6500 1817 6556
rect 1817 6500 1821 6556
rect 1757 6496 1821 6500
rect 1837 6556 1901 6560
rect 1837 6500 1841 6556
rect 1841 6500 1897 6556
rect 1897 6500 1901 6556
rect 1837 6496 1901 6500
rect 1917 6556 1981 6560
rect 1917 6500 1921 6556
rect 1921 6500 1977 6556
rect 1977 6500 1981 6556
rect 1917 6496 1981 6500
rect 1997 6556 2061 6560
rect 1997 6500 2001 6556
rect 2001 6500 2057 6556
rect 2057 6500 2061 6556
rect 1997 6496 2061 6500
rect 4471 6556 4535 6560
rect 4471 6500 4475 6556
rect 4475 6500 4531 6556
rect 4531 6500 4535 6556
rect 4471 6496 4535 6500
rect 4551 6556 4615 6560
rect 4551 6500 4555 6556
rect 4555 6500 4611 6556
rect 4611 6500 4615 6556
rect 4551 6496 4615 6500
rect 4631 6556 4695 6560
rect 4631 6500 4635 6556
rect 4635 6500 4691 6556
rect 4691 6500 4695 6556
rect 4631 6496 4695 6500
rect 4711 6556 4775 6560
rect 4711 6500 4715 6556
rect 4715 6500 4771 6556
rect 4771 6500 4775 6556
rect 4711 6496 4775 6500
rect 7185 6556 7249 6560
rect 7185 6500 7189 6556
rect 7189 6500 7245 6556
rect 7245 6500 7249 6556
rect 7185 6496 7249 6500
rect 7265 6556 7329 6560
rect 7265 6500 7269 6556
rect 7269 6500 7325 6556
rect 7325 6500 7329 6556
rect 7265 6496 7329 6500
rect 7345 6556 7409 6560
rect 7345 6500 7349 6556
rect 7349 6500 7405 6556
rect 7405 6500 7409 6556
rect 7345 6496 7409 6500
rect 7425 6556 7489 6560
rect 7425 6500 7429 6556
rect 7429 6500 7485 6556
rect 7485 6500 7489 6556
rect 7425 6496 7489 6500
rect 9899 6556 9963 6560
rect 9899 6500 9903 6556
rect 9903 6500 9959 6556
rect 9959 6500 9963 6556
rect 9899 6496 9963 6500
rect 9979 6556 10043 6560
rect 9979 6500 9983 6556
rect 9983 6500 10039 6556
rect 10039 6500 10043 6556
rect 9979 6496 10043 6500
rect 10059 6556 10123 6560
rect 10059 6500 10063 6556
rect 10063 6500 10119 6556
rect 10119 6500 10123 6556
rect 10059 6496 10123 6500
rect 10139 6556 10203 6560
rect 10139 6500 10143 6556
rect 10143 6500 10199 6556
rect 10199 6500 10203 6556
rect 10139 6496 10203 6500
rect 7604 6080 7668 6084
rect 7604 6024 7618 6080
rect 7618 6024 7668 6080
rect 7604 6020 7668 6024
rect 3114 6012 3178 6016
rect 3114 5956 3118 6012
rect 3118 5956 3174 6012
rect 3174 5956 3178 6012
rect 3114 5952 3178 5956
rect 3194 6012 3258 6016
rect 3194 5956 3198 6012
rect 3198 5956 3254 6012
rect 3254 5956 3258 6012
rect 3194 5952 3258 5956
rect 3274 6012 3338 6016
rect 3274 5956 3278 6012
rect 3278 5956 3334 6012
rect 3334 5956 3338 6012
rect 3274 5952 3338 5956
rect 3354 6012 3418 6016
rect 3354 5956 3358 6012
rect 3358 5956 3414 6012
rect 3414 5956 3418 6012
rect 3354 5952 3418 5956
rect 5828 6012 5892 6016
rect 5828 5956 5832 6012
rect 5832 5956 5888 6012
rect 5888 5956 5892 6012
rect 5828 5952 5892 5956
rect 5908 6012 5972 6016
rect 5908 5956 5912 6012
rect 5912 5956 5968 6012
rect 5968 5956 5972 6012
rect 5908 5952 5972 5956
rect 5988 6012 6052 6016
rect 5988 5956 5992 6012
rect 5992 5956 6048 6012
rect 6048 5956 6052 6012
rect 5988 5952 6052 5956
rect 6068 6012 6132 6016
rect 6068 5956 6072 6012
rect 6072 5956 6128 6012
rect 6128 5956 6132 6012
rect 6068 5952 6132 5956
rect 8542 6012 8606 6016
rect 8542 5956 8546 6012
rect 8546 5956 8602 6012
rect 8602 5956 8606 6012
rect 8542 5952 8606 5956
rect 8622 6012 8686 6016
rect 8622 5956 8626 6012
rect 8626 5956 8682 6012
rect 8682 5956 8686 6012
rect 8622 5952 8686 5956
rect 8702 6012 8766 6016
rect 8702 5956 8706 6012
rect 8706 5956 8762 6012
rect 8762 5956 8766 6012
rect 8702 5952 8766 5956
rect 8782 6012 8846 6016
rect 8782 5956 8786 6012
rect 8786 5956 8842 6012
rect 8842 5956 8846 6012
rect 8782 5952 8846 5956
rect 11256 6012 11320 6016
rect 11256 5956 11260 6012
rect 11260 5956 11316 6012
rect 11316 5956 11320 6012
rect 11256 5952 11320 5956
rect 11336 6012 11400 6016
rect 11336 5956 11340 6012
rect 11340 5956 11396 6012
rect 11396 5956 11400 6012
rect 11336 5952 11400 5956
rect 11416 6012 11480 6016
rect 11416 5956 11420 6012
rect 11420 5956 11476 6012
rect 11476 5956 11480 6012
rect 11416 5952 11480 5956
rect 11496 6012 11560 6016
rect 11496 5956 11500 6012
rect 11500 5956 11556 6012
rect 11556 5956 11560 6012
rect 11496 5952 11560 5956
rect 1757 5468 1821 5472
rect 1757 5412 1761 5468
rect 1761 5412 1817 5468
rect 1817 5412 1821 5468
rect 1757 5408 1821 5412
rect 1837 5468 1901 5472
rect 1837 5412 1841 5468
rect 1841 5412 1897 5468
rect 1897 5412 1901 5468
rect 1837 5408 1901 5412
rect 1917 5468 1981 5472
rect 1917 5412 1921 5468
rect 1921 5412 1977 5468
rect 1977 5412 1981 5468
rect 1917 5408 1981 5412
rect 1997 5468 2061 5472
rect 1997 5412 2001 5468
rect 2001 5412 2057 5468
rect 2057 5412 2061 5468
rect 1997 5408 2061 5412
rect 4471 5468 4535 5472
rect 4471 5412 4475 5468
rect 4475 5412 4531 5468
rect 4531 5412 4535 5468
rect 4471 5408 4535 5412
rect 4551 5468 4615 5472
rect 4551 5412 4555 5468
rect 4555 5412 4611 5468
rect 4611 5412 4615 5468
rect 4551 5408 4615 5412
rect 4631 5468 4695 5472
rect 4631 5412 4635 5468
rect 4635 5412 4691 5468
rect 4691 5412 4695 5468
rect 4631 5408 4695 5412
rect 4711 5468 4775 5472
rect 4711 5412 4715 5468
rect 4715 5412 4771 5468
rect 4771 5412 4775 5468
rect 4711 5408 4775 5412
rect 7185 5468 7249 5472
rect 7185 5412 7189 5468
rect 7189 5412 7245 5468
rect 7245 5412 7249 5468
rect 7185 5408 7249 5412
rect 7265 5468 7329 5472
rect 7265 5412 7269 5468
rect 7269 5412 7325 5468
rect 7325 5412 7329 5468
rect 7265 5408 7329 5412
rect 7345 5468 7409 5472
rect 7345 5412 7349 5468
rect 7349 5412 7405 5468
rect 7405 5412 7409 5468
rect 7345 5408 7409 5412
rect 7425 5468 7489 5472
rect 7425 5412 7429 5468
rect 7429 5412 7485 5468
rect 7485 5412 7489 5468
rect 7425 5408 7489 5412
rect 9899 5468 9963 5472
rect 9899 5412 9903 5468
rect 9903 5412 9959 5468
rect 9959 5412 9963 5468
rect 9899 5408 9963 5412
rect 9979 5468 10043 5472
rect 9979 5412 9983 5468
rect 9983 5412 10039 5468
rect 10039 5412 10043 5468
rect 9979 5408 10043 5412
rect 10059 5468 10123 5472
rect 10059 5412 10063 5468
rect 10063 5412 10119 5468
rect 10119 5412 10123 5468
rect 10059 5408 10123 5412
rect 10139 5468 10203 5472
rect 10139 5412 10143 5468
rect 10143 5412 10199 5468
rect 10199 5412 10203 5468
rect 10139 5408 10203 5412
rect 3114 4924 3178 4928
rect 3114 4868 3118 4924
rect 3118 4868 3174 4924
rect 3174 4868 3178 4924
rect 3114 4864 3178 4868
rect 3194 4924 3258 4928
rect 3194 4868 3198 4924
rect 3198 4868 3254 4924
rect 3254 4868 3258 4924
rect 3194 4864 3258 4868
rect 3274 4924 3338 4928
rect 3274 4868 3278 4924
rect 3278 4868 3334 4924
rect 3334 4868 3338 4924
rect 3274 4864 3338 4868
rect 3354 4924 3418 4928
rect 3354 4868 3358 4924
rect 3358 4868 3414 4924
rect 3414 4868 3418 4924
rect 3354 4864 3418 4868
rect 5828 4924 5892 4928
rect 5828 4868 5832 4924
rect 5832 4868 5888 4924
rect 5888 4868 5892 4924
rect 5828 4864 5892 4868
rect 5908 4924 5972 4928
rect 5908 4868 5912 4924
rect 5912 4868 5968 4924
rect 5968 4868 5972 4924
rect 5908 4864 5972 4868
rect 5988 4924 6052 4928
rect 5988 4868 5992 4924
rect 5992 4868 6048 4924
rect 6048 4868 6052 4924
rect 5988 4864 6052 4868
rect 6068 4924 6132 4928
rect 6068 4868 6072 4924
rect 6072 4868 6128 4924
rect 6128 4868 6132 4924
rect 6068 4864 6132 4868
rect 8542 4924 8606 4928
rect 8542 4868 8546 4924
rect 8546 4868 8602 4924
rect 8602 4868 8606 4924
rect 8542 4864 8606 4868
rect 8622 4924 8686 4928
rect 8622 4868 8626 4924
rect 8626 4868 8682 4924
rect 8682 4868 8686 4924
rect 8622 4864 8686 4868
rect 8702 4924 8766 4928
rect 8702 4868 8706 4924
rect 8706 4868 8762 4924
rect 8762 4868 8766 4924
rect 8702 4864 8766 4868
rect 8782 4924 8846 4928
rect 8782 4868 8786 4924
rect 8786 4868 8842 4924
rect 8842 4868 8846 4924
rect 8782 4864 8846 4868
rect 11256 4924 11320 4928
rect 11256 4868 11260 4924
rect 11260 4868 11316 4924
rect 11316 4868 11320 4924
rect 11256 4864 11320 4868
rect 11336 4924 11400 4928
rect 11336 4868 11340 4924
rect 11340 4868 11396 4924
rect 11396 4868 11400 4924
rect 11336 4864 11400 4868
rect 11416 4924 11480 4928
rect 11416 4868 11420 4924
rect 11420 4868 11476 4924
rect 11476 4868 11480 4924
rect 11416 4864 11480 4868
rect 11496 4924 11560 4928
rect 11496 4868 11500 4924
rect 11500 4868 11556 4924
rect 11556 4868 11560 4924
rect 11496 4864 11560 4868
rect 1757 4380 1821 4384
rect 1757 4324 1761 4380
rect 1761 4324 1817 4380
rect 1817 4324 1821 4380
rect 1757 4320 1821 4324
rect 1837 4380 1901 4384
rect 1837 4324 1841 4380
rect 1841 4324 1897 4380
rect 1897 4324 1901 4380
rect 1837 4320 1901 4324
rect 1917 4380 1981 4384
rect 1917 4324 1921 4380
rect 1921 4324 1977 4380
rect 1977 4324 1981 4380
rect 1917 4320 1981 4324
rect 1997 4380 2061 4384
rect 1997 4324 2001 4380
rect 2001 4324 2057 4380
rect 2057 4324 2061 4380
rect 1997 4320 2061 4324
rect 4471 4380 4535 4384
rect 4471 4324 4475 4380
rect 4475 4324 4531 4380
rect 4531 4324 4535 4380
rect 4471 4320 4535 4324
rect 4551 4380 4615 4384
rect 4551 4324 4555 4380
rect 4555 4324 4611 4380
rect 4611 4324 4615 4380
rect 4551 4320 4615 4324
rect 4631 4380 4695 4384
rect 4631 4324 4635 4380
rect 4635 4324 4691 4380
rect 4691 4324 4695 4380
rect 4631 4320 4695 4324
rect 4711 4380 4775 4384
rect 4711 4324 4715 4380
rect 4715 4324 4771 4380
rect 4771 4324 4775 4380
rect 4711 4320 4775 4324
rect 7185 4380 7249 4384
rect 7185 4324 7189 4380
rect 7189 4324 7245 4380
rect 7245 4324 7249 4380
rect 7185 4320 7249 4324
rect 7265 4380 7329 4384
rect 7265 4324 7269 4380
rect 7269 4324 7325 4380
rect 7325 4324 7329 4380
rect 7265 4320 7329 4324
rect 7345 4380 7409 4384
rect 7345 4324 7349 4380
rect 7349 4324 7405 4380
rect 7405 4324 7409 4380
rect 7345 4320 7409 4324
rect 7425 4380 7489 4384
rect 7425 4324 7429 4380
rect 7429 4324 7485 4380
rect 7485 4324 7489 4380
rect 7425 4320 7489 4324
rect 9899 4380 9963 4384
rect 9899 4324 9903 4380
rect 9903 4324 9959 4380
rect 9959 4324 9963 4380
rect 9899 4320 9963 4324
rect 9979 4380 10043 4384
rect 9979 4324 9983 4380
rect 9983 4324 10039 4380
rect 10039 4324 10043 4380
rect 9979 4320 10043 4324
rect 10059 4380 10123 4384
rect 10059 4324 10063 4380
rect 10063 4324 10119 4380
rect 10119 4324 10123 4380
rect 10059 4320 10123 4324
rect 10139 4380 10203 4384
rect 10139 4324 10143 4380
rect 10143 4324 10199 4380
rect 10199 4324 10203 4380
rect 10139 4320 10203 4324
rect 3114 3836 3178 3840
rect 3114 3780 3118 3836
rect 3118 3780 3174 3836
rect 3174 3780 3178 3836
rect 3114 3776 3178 3780
rect 3194 3836 3258 3840
rect 3194 3780 3198 3836
rect 3198 3780 3254 3836
rect 3254 3780 3258 3836
rect 3194 3776 3258 3780
rect 3274 3836 3338 3840
rect 3274 3780 3278 3836
rect 3278 3780 3334 3836
rect 3334 3780 3338 3836
rect 3274 3776 3338 3780
rect 3354 3836 3418 3840
rect 3354 3780 3358 3836
rect 3358 3780 3414 3836
rect 3414 3780 3418 3836
rect 3354 3776 3418 3780
rect 5828 3836 5892 3840
rect 5828 3780 5832 3836
rect 5832 3780 5888 3836
rect 5888 3780 5892 3836
rect 5828 3776 5892 3780
rect 5908 3836 5972 3840
rect 5908 3780 5912 3836
rect 5912 3780 5968 3836
rect 5968 3780 5972 3836
rect 5908 3776 5972 3780
rect 5988 3836 6052 3840
rect 5988 3780 5992 3836
rect 5992 3780 6048 3836
rect 6048 3780 6052 3836
rect 5988 3776 6052 3780
rect 6068 3836 6132 3840
rect 6068 3780 6072 3836
rect 6072 3780 6128 3836
rect 6128 3780 6132 3836
rect 6068 3776 6132 3780
rect 8542 3836 8606 3840
rect 8542 3780 8546 3836
rect 8546 3780 8602 3836
rect 8602 3780 8606 3836
rect 8542 3776 8606 3780
rect 8622 3836 8686 3840
rect 8622 3780 8626 3836
rect 8626 3780 8682 3836
rect 8682 3780 8686 3836
rect 8622 3776 8686 3780
rect 8702 3836 8766 3840
rect 8702 3780 8706 3836
rect 8706 3780 8762 3836
rect 8762 3780 8766 3836
rect 8702 3776 8766 3780
rect 8782 3836 8846 3840
rect 8782 3780 8786 3836
rect 8786 3780 8842 3836
rect 8842 3780 8846 3836
rect 8782 3776 8846 3780
rect 11256 3836 11320 3840
rect 11256 3780 11260 3836
rect 11260 3780 11316 3836
rect 11316 3780 11320 3836
rect 11256 3776 11320 3780
rect 11336 3836 11400 3840
rect 11336 3780 11340 3836
rect 11340 3780 11396 3836
rect 11396 3780 11400 3836
rect 11336 3776 11400 3780
rect 11416 3836 11480 3840
rect 11416 3780 11420 3836
rect 11420 3780 11476 3836
rect 11476 3780 11480 3836
rect 11416 3776 11480 3780
rect 11496 3836 11560 3840
rect 11496 3780 11500 3836
rect 11500 3780 11556 3836
rect 11556 3780 11560 3836
rect 11496 3776 11560 3780
rect 1757 3292 1821 3296
rect 1757 3236 1761 3292
rect 1761 3236 1817 3292
rect 1817 3236 1821 3292
rect 1757 3232 1821 3236
rect 1837 3292 1901 3296
rect 1837 3236 1841 3292
rect 1841 3236 1897 3292
rect 1897 3236 1901 3292
rect 1837 3232 1901 3236
rect 1917 3292 1981 3296
rect 1917 3236 1921 3292
rect 1921 3236 1977 3292
rect 1977 3236 1981 3292
rect 1917 3232 1981 3236
rect 1997 3292 2061 3296
rect 1997 3236 2001 3292
rect 2001 3236 2057 3292
rect 2057 3236 2061 3292
rect 1997 3232 2061 3236
rect 4471 3292 4535 3296
rect 4471 3236 4475 3292
rect 4475 3236 4531 3292
rect 4531 3236 4535 3292
rect 4471 3232 4535 3236
rect 4551 3292 4615 3296
rect 4551 3236 4555 3292
rect 4555 3236 4611 3292
rect 4611 3236 4615 3292
rect 4551 3232 4615 3236
rect 4631 3292 4695 3296
rect 4631 3236 4635 3292
rect 4635 3236 4691 3292
rect 4691 3236 4695 3292
rect 4631 3232 4695 3236
rect 4711 3292 4775 3296
rect 4711 3236 4715 3292
rect 4715 3236 4771 3292
rect 4771 3236 4775 3292
rect 4711 3232 4775 3236
rect 7185 3292 7249 3296
rect 7185 3236 7189 3292
rect 7189 3236 7245 3292
rect 7245 3236 7249 3292
rect 7185 3232 7249 3236
rect 7265 3292 7329 3296
rect 7265 3236 7269 3292
rect 7269 3236 7325 3292
rect 7325 3236 7329 3292
rect 7265 3232 7329 3236
rect 7345 3292 7409 3296
rect 7345 3236 7349 3292
rect 7349 3236 7405 3292
rect 7405 3236 7409 3292
rect 7345 3232 7409 3236
rect 7425 3292 7489 3296
rect 7425 3236 7429 3292
rect 7429 3236 7485 3292
rect 7485 3236 7489 3292
rect 7425 3232 7489 3236
rect 9899 3292 9963 3296
rect 9899 3236 9903 3292
rect 9903 3236 9959 3292
rect 9959 3236 9963 3292
rect 9899 3232 9963 3236
rect 9979 3292 10043 3296
rect 9979 3236 9983 3292
rect 9983 3236 10039 3292
rect 10039 3236 10043 3292
rect 9979 3232 10043 3236
rect 10059 3292 10123 3296
rect 10059 3236 10063 3292
rect 10063 3236 10119 3292
rect 10119 3236 10123 3292
rect 10059 3232 10123 3236
rect 10139 3292 10203 3296
rect 10139 3236 10143 3292
rect 10143 3236 10199 3292
rect 10199 3236 10203 3292
rect 10139 3232 10203 3236
rect 3114 2748 3178 2752
rect 3114 2692 3118 2748
rect 3118 2692 3174 2748
rect 3174 2692 3178 2748
rect 3114 2688 3178 2692
rect 3194 2748 3258 2752
rect 3194 2692 3198 2748
rect 3198 2692 3254 2748
rect 3254 2692 3258 2748
rect 3194 2688 3258 2692
rect 3274 2748 3338 2752
rect 3274 2692 3278 2748
rect 3278 2692 3334 2748
rect 3334 2692 3338 2748
rect 3274 2688 3338 2692
rect 3354 2748 3418 2752
rect 3354 2692 3358 2748
rect 3358 2692 3414 2748
rect 3414 2692 3418 2748
rect 3354 2688 3418 2692
rect 5828 2748 5892 2752
rect 5828 2692 5832 2748
rect 5832 2692 5888 2748
rect 5888 2692 5892 2748
rect 5828 2688 5892 2692
rect 5908 2748 5972 2752
rect 5908 2692 5912 2748
rect 5912 2692 5968 2748
rect 5968 2692 5972 2748
rect 5908 2688 5972 2692
rect 5988 2748 6052 2752
rect 5988 2692 5992 2748
rect 5992 2692 6048 2748
rect 6048 2692 6052 2748
rect 5988 2688 6052 2692
rect 6068 2748 6132 2752
rect 6068 2692 6072 2748
rect 6072 2692 6128 2748
rect 6128 2692 6132 2748
rect 6068 2688 6132 2692
rect 8542 2748 8606 2752
rect 8542 2692 8546 2748
rect 8546 2692 8602 2748
rect 8602 2692 8606 2748
rect 8542 2688 8606 2692
rect 8622 2748 8686 2752
rect 8622 2692 8626 2748
rect 8626 2692 8682 2748
rect 8682 2692 8686 2748
rect 8622 2688 8686 2692
rect 8702 2748 8766 2752
rect 8702 2692 8706 2748
rect 8706 2692 8762 2748
rect 8762 2692 8766 2748
rect 8702 2688 8766 2692
rect 8782 2748 8846 2752
rect 8782 2692 8786 2748
rect 8786 2692 8842 2748
rect 8842 2692 8846 2748
rect 8782 2688 8846 2692
rect 11256 2748 11320 2752
rect 11256 2692 11260 2748
rect 11260 2692 11316 2748
rect 11316 2692 11320 2748
rect 11256 2688 11320 2692
rect 11336 2748 11400 2752
rect 11336 2692 11340 2748
rect 11340 2692 11396 2748
rect 11396 2692 11400 2748
rect 11336 2688 11400 2692
rect 11416 2748 11480 2752
rect 11416 2692 11420 2748
rect 11420 2692 11476 2748
rect 11476 2692 11480 2748
rect 11416 2688 11480 2692
rect 11496 2748 11560 2752
rect 11496 2692 11500 2748
rect 11500 2692 11556 2748
rect 11556 2692 11560 2748
rect 11496 2688 11560 2692
rect 7604 2484 7668 2548
rect 1757 2204 1821 2208
rect 1757 2148 1761 2204
rect 1761 2148 1817 2204
rect 1817 2148 1821 2204
rect 1757 2144 1821 2148
rect 1837 2204 1901 2208
rect 1837 2148 1841 2204
rect 1841 2148 1897 2204
rect 1897 2148 1901 2204
rect 1837 2144 1901 2148
rect 1917 2204 1981 2208
rect 1917 2148 1921 2204
rect 1921 2148 1977 2204
rect 1977 2148 1981 2204
rect 1917 2144 1981 2148
rect 1997 2204 2061 2208
rect 1997 2148 2001 2204
rect 2001 2148 2057 2204
rect 2057 2148 2061 2204
rect 1997 2144 2061 2148
rect 4471 2204 4535 2208
rect 4471 2148 4475 2204
rect 4475 2148 4531 2204
rect 4531 2148 4535 2204
rect 4471 2144 4535 2148
rect 4551 2204 4615 2208
rect 4551 2148 4555 2204
rect 4555 2148 4611 2204
rect 4611 2148 4615 2204
rect 4551 2144 4615 2148
rect 4631 2204 4695 2208
rect 4631 2148 4635 2204
rect 4635 2148 4691 2204
rect 4691 2148 4695 2204
rect 4631 2144 4695 2148
rect 4711 2204 4775 2208
rect 4711 2148 4715 2204
rect 4715 2148 4771 2204
rect 4771 2148 4775 2204
rect 4711 2144 4775 2148
rect 7185 2204 7249 2208
rect 7185 2148 7189 2204
rect 7189 2148 7245 2204
rect 7245 2148 7249 2204
rect 7185 2144 7249 2148
rect 7265 2204 7329 2208
rect 7265 2148 7269 2204
rect 7269 2148 7325 2204
rect 7325 2148 7329 2204
rect 7265 2144 7329 2148
rect 7345 2204 7409 2208
rect 7345 2148 7349 2204
rect 7349 2148 7405 2204
rect 7405 2148 7409 2204
rect 7345 2144 7409 2148
rect 7425 2204 7489 2208
rect 7425 2148 7429 2204
rect 7429 2148 7485 2204
rect 7485 2148 7489 2204
rect 7425 2144 7489 2148
rect 9899 2204 9963 2208
rect 9899 2148 9903 2204
rect 9903 2148 9959 2204
rect 9959 2148 9963 2204
rect 9899 2144 9963 2148
rect 9979 2204 10043 2208
rect 9979 2148 9983 2204
rect 9983 2148 10039 2204
rect 10039 2148 10043 2204
rect 9979 2144 10043 2148
rect 10059 2204 10123 2208
rect 10059 2148 10063 2204
rect 10063 2148 10119 2204
rect 10119 2148 10123 2204
rect 10059 2144 10123 2148
rect 10139 2204 10203 2208
rect 10139 2148 10143 2204
rect 10143 2148 10199 2204
rect 10199 2148 10203 2204
rect 10139 2144 10203 2148
rect 3114 1660 3178 1664
rect 3114 1604 3118 1660
rect 3118 1604 3174 1660
rect 3174 1604 3178 1660
rect 3114 1600 3178 1604
rect 3194 1660 3258 1664
rect 3194 1604 3198 1660
rect 3198 1604 3254 1660
rect 3254 1604 3258 1660
rect 3194 1600 3258 1604
rect 3274 1660 3338 1664
rect 3274 1604 3278 1660
rect 3278 1604 3334 1660
rect 3334 1604 3338 1660
rect 3274 1600 3338 1604
rect 3354 1660 3418 1664
rect 3354 1604 3358 1660
rect 3358 1604 3414 1660
rect 3414 1604 3418 1660
rect 3354 1600 3418 1604
rect 5828 1660 5892 1664
rect 5828 1604 5832 1660
rect 5832 1604 5888 1660
rect 5888 1604 5892 1660
rect 5828 1600 5892 1604
rect 5908 1660 5972 1664
rect 5908 1604 5912 1660
rect 5912 1604 5968 1660
rect 5968 1604 5972 1660
rect 5908 1600 5972 1604
rect 5988 1660 6052 1664
rect 5988 1604 5992 1660
rect 5992 1604 6048 1660
rect 6048 1604 6052 1660
rect 5988 1600 6052 1604
rect 6068 1660 6132 1664
rect 6068 1604 6072 1660
rect 6072 1604 6128 1660
rect 6128 1604 6132 1660
rect 6068 1600 6132 1604
rect 8542 1660 8606 1664
rect 8542 1604 8546 1660
rect 8546 1604 8602 1660
rect 8602 1604 8606 1660
rect 8542 1600 8606 1604
rect 8622 1660 8686 1664
rect 8622 1604 8626 1660
rect 8626 1604 8682 1660
rect 8682 1604 8686 1660
rect 8622 1600 8686 1604
rect 8702 1660 8766 1664
rect 8702 1604 8706 1660
rect 8706 1604 8762 1660
rect 8762 1604 8766 1660
rect 8702 1600 8766 1604
rect 8782 1660 8846 1664
rect 8782 1604 8786 1660
rect 8786 1604 8842 1660
rect 8842 1604 8846 1660
rect 8782 1600 8846 1604
rect 11256 1660 11320 1664
rect 11256 1604 11260 1660
rect 11260 1604 11316 1660
rect 11316 1604 11320 1660
rect 11256 1600 11320 1604
rect 11336 1660 11400 1664
rect 11336 1604 11340 1660
rect 11340 1604 11396 1660
rect 11396 1604 11400 1660
rect 11336 1600 11400 1604
rect 11416 1660 11480 1664
rect 11416 1604 11420 1660
rect 11420 1604 11476 1660
rect 11476 1604 11480 1660
rect 11416 1600 11480 1604
rect 11496 1660 11560 1664
rect 11496 1604 11500 1660
rect 11500 1604 11556 1660
rect 11556 1604 11560 1660
rect 11496 1600 11560 1604
rect 1757 1116 1821 1120
rect 1757 1060 1761 1116
rect 1761 1060 1817 1116
rect 1817 1060 1821 1116
rect 1757 1056 1821 1060
rect 1837 1116 1901 1120
rect 1837 1060 1841 1116
rect 1841 1060 1897 1116
rect 1897 1060 1901 1116
rect 1837 1056 1901 1060
rect 1917 1116 1981 1120
rect 1917 1060 1921 1116
rect 1921 1060 1977 1116
rect 1977 1060 1981 1116
rect 1917 1056 1981 1060
rect 1997 1116 2061 1120
rect 1997 1060 2001 1116
rect 2001 1060 2057 1116
rect 2057 1060 2061 1116
rect 1997 1056 2061 1060
rect 4471 1116 4535 1120
rect 4471 1060 4475 1116
rect 4475 1060 4531 1116
rect 4531 1060 4535 1116
rect 4471 1056 4535 1060
rect 4551 1116 4615 1120
rect 4551 1060 4555 1116
rect 4555 1060 4611 1116
rect 4611 1060 4615 1116
rect 4551 1056 4615 1060
rect 4631 1116 4695 1120
rect 4631 1060 4635 1116
rect 4635 1060 4691 1116
rect 4691 1060 4695 1116
rect 4631 1056 4695 1060
rect 4711 1116 4775 1120
rect 4711 1060 4715 1116
rect 4715 1060 4771 1116
rect 4771 1060 4775 1116
rect 4711 1056 4775 1060
rect 7185 1116 7249 1120
rect 7185 1060 7189 1116
rect 7189 1060 7245 1116
rect 7245 1060 7249 1116
rect 7185 1056 7249 1060
rect 7265 1116 7329 1120
rect 7265 1060 7269 1116
rect 7269 1060 7325 1116
rect 7325 1060 7329 1116
rect 7265 1056 7329 1060
rect 7345 1116 7409 1120
rect 7345 1060 7349 1116
rect 7349 1060 7405 1116
rect 7405 1060 7409 1116
rect 7345 1056 7409 1060
rect 7425 1116 7489 1120
rect 7425 1060 7429 1116
rect 7429 1060 7485 1116
rect 7485 1060 7489 1116
rect 7425 1056 7489 1060
rect 9899 1116 9963 1120
rect 9899 1060 9903 1116
rect 9903 1060 9959 1116
rect 9959 1060 9963 1116
rect 9899 1056 9963 1060
rect 9979 1116 10043 1120
rect 9979 1060 9983 1116
rect 9983 1060 10039 1116
rect 10039 1060 10043 1116
rect 9979 1056 10043 1060
rect 10059 1116 10123 1120
rect 10059 1060 10063 1116
rect 10063 1060 10119 1116
rect 10119 1060 10123 1116
rect 10059 1056 10123 1060
rect 10139 1116 10203 1120
rect 10139 1060 10143 1116
rect 10143 1060 10199 1116
rect 10199 1060 10203 1116
rect 10139 1056 10203 1060
rect 3114 572 3178 576
rect 3114 516 3118 572
rect 3118 516 3174 572
rect 3174 516 3178 572
rect 3114 512 3178 516
rect 3194 572 3258 576
rect 3194 516 3198 572
rect 3198 516 3254 572
rect 3254 516 3258 572
rect 3194 512 3258 516
rect 3274 572 3338 576
rect 3274 516 3278 572
rect 3278 516 3334 572
rect 3334 516 3338 572
rect 3274 512 3338 516
rect 3354 572 3418 576
rect 3354 516 3358 572
rect 3358 516 3414 572
rect 3414 516 3418 572
rect 3354 512 3418 516
rect 5828 572 5892 576
rect 5828 516 5832 572
rect 5832 516 5888 572
rect 5888 516 5892 572
rect 5828 512 5892 516
rect 5908 572 5972 576
rect 5908 516 5912 572
rect 5912 516 5968 572
rect 5968 516 5972 572
rect 5908 512 5972 516
rect 5988 572 6052 576
rect 5988 516 5992 572
rect 5992 516 6048 572
rect 6048 516 6052 572
rect 5988 512 6052 516
rect 6068 572 6132 576
rect 6068 516 6072 572
rect 6072 516 6128 572
rect 6128 516 6132 572
rect 6068 512 6132 516
rect 8542 572 8606 576
rect 8542 516 8546 572
rect 8546 516 8602 572
rect 8602 516 8606 572
rect 8542 512 8606 516
rect 8622 572 8686 576
rect 8622 516 8626 572
rect 8626 516 8682 572
rect 8682 516 8686 572
rect 8622 512 8686 516
rect 8702 572 8766 576
rect 8702 516 8706 572
rect 8706 516 8762 572
rect 8762 516 8766 572
rect 8702 512 8766 516
rect 8782 572 8846 576
rect 8782 516 8786 572
rect 8786 516 8842 572
rect 8842 516 8846 572
rect 8782 512 8846 516
rect 11256 572 11320 576
rect 11256 516 11260 572
rect 11260 516 11316 572
rect 11316 516 11320 572
rect 11256 512 11320 516
rect 11336 572 11400 576
rect 11336 516 11340 572
rect 11340 516 11396 572
rect 11396 516 11400 572
rect 11336 512 11400 516
rect 11416 572 11480 576
rect 11416 516 11420 572
rect 11420 516 11476 572
rect 11476 516 11480 572
rect 11416 512 11480 516
rect 11496 572 11560 576
rect 11496 516 11500 572
rect 11500 516 11556 572
rect 11556 516 11560 572
rect 11496 512 11560 516
<< metal4 >>
rect 1749 8736 2069 9296
rect 1749 8672 1757 8736
rect 1821 8672 1837 8736
rect 1901 8672 1917 8736
rect 1981 8672 1997 8736
rect 2061 8672 2069 8736
rect 1749 7648 2069 8672
rect 1749 7584 1757 7648
rect 1821 7584 1837 7648
rect 1901 7584 1917 7648
rect 1981 7584 1997 7648
rect 2061 7584 2069 7648
rect 1749 6560 2069 7584
rect 1749 6496 1757 6560
rect 1821 6496 1837 6560
rect 1901 6496 1917 6560
rect 1981 6496 1997 6560
rect 2061 6496 2069 6560
rect 1749 5472 2069 6496
rect 1749 5408 1757 5472
rect 1821 5408 1837 5472
rect 1901 5408 1917 5472
rect 1981 5408 1997 5472
rect 2061 5408 2069 5472
rect 1749 4384 2069 5408
rect 1749 4320 1757 4384
rect 1821 4320 1837 4384
rect 1901 4320 1917 4384
rect 1981 4320 1997 4384
rect 2061 4320 2069 4384
rect 1749 3296 2069 4320
rect 1749 3232 1757 3296
rect 1821 3232 1837 3296
rect 1901 3232 1917 3296
rect 1981 3232 1997 3296
rect 2061 3232 2069 3296
rect 1749 2208 2069 3232
rect 1749 2144 1757 2208
rect 1821 2144 1837 2208
rect 1901 2144 1917 2208
rect 1981 2144 1997 2208
rect 2061 2144 2069 2208
rect 1749 1120 2069 2144
rect 1749 1056 1757 1120
rect 1821 1056 1837 1120
rect 1901 1056 1917 1120
rect 1981 1056 1997 1120
rect 2061 1056 2069 1120
rect 1749 496 2069 1056
rect 3106 9280 3426 9296
rect 3106 9216 3114 9280
rect 3178 9216 3194 9280
rect 3258 9216 3274 9280
rect 3338 9216 3354 9280
rect 3418 9216 3426 9280
rect 3106 8192 3426 9216
rect 3106 8128 3114 8192
rect 3178 8128 3194 8192
rect 3258 8128 3274 8192
rect 3338 8128 3354 8192
rect 3418 8128 3426 8192
rect 3106 7104 3426 8128
rect 3106 7040 3114 7104
rect 3178 7040 3194 7104
rect 3258 7040 3274 7104
rect 3338 7040 3354 7104
rect 3418 7040 3426 7104
rect 3106 6016 3426 7040
rect 3106 5952 3114 6016
rect 3178 5952 3194 6016
rect 3258 5952 3274 6016
rect 3338 5952 3354 6016
rect 3418 5952 3426 6016
rect 3106 4928 3426 5952
rect 3106 4864 3114 4928
rect 3178 4864 3194 4928
rect 3258 4864 3274 4928
rect 3338 4864 3354 4928
rect 3418 4864 3426 4928
rect 3106 3840 3426 4864
rect 3106 3776 3114 3840
rect 3178 3776 3194 3840
rect 3258 3776 3274 3840
rect 3338 3776 3354 3840
rect 3418 3776 3426 3840
rect 3106 2752 3426 3776
rect 3106 2688 3114 2752
rect 3178 2688 3194 2752
rect 3258 2688 3274 2752
rect 3338 2688 3354 2752
rect 3418 2688 3426 2752
rect 3106 1664 3426 2688
rect 3106 1600 3114 1664
rect 3178 1600 3194 1664
rect 3258 1600 3274 1664
rect 3338 1600 3354 1664
rect 3418 1600 3426 1664
rect 3106 576 3426 1600
rect 3106 512 3114 576
rect 3178 512 3194 576
rect 3258 512 3274 576
rect 3338 512 3354 576
rect 3418 512 3426 576
rect 3106 496 3426 512
rect 4463 8736 4783 9296
rect 4463 8672 4471 8736
rect 4535 8672 4551 8736
rect 4615 8672 4631 8736
rect 4695 8672 4711 8736
rect 4775 8672 4783 8736
rect 4463 7648 4783 8672
rect 4463 7584 4471 7648
rect 4535 7584 4551 7648
rect 4615 7584 4631 7648
rect 4695 7584 4711 7648
rect 4775 7584 4783 7648
rect 4463 6560 4783 7584
rect 4463 6496 4471 6560
rect 4535 6496 4551 6560
rect 4615 6496 4631 6560
rect 4695 6496 4711 6560
rect 4775 6496 4783 6560
rect 4463 5472 4783 6496
rect 4463 5408 4471 5472
rect 4535 5408 4551 5472
rect 4615 5408 4631 5472
rect 4695 5408 4711 5472
rect 4775 5408 4783 5472
rect 4463 4384 4783 5408
rect 4463 4320 4471 4384
rect 4535 4320 4551 4384
rect 4615 4320 4631 4384
rect 4695 4320 4711 4384
rect 4775 4320 4783 4384
rect 4463 3296 4783 4320
rect 4463 3232 4471 3296
rect 4535 3232 4551 3296
rect 4615 3232 4631 3296
rect 4695 3232 4711 3296
rect 4775 3232 4783 3296
rect 4463 2208 4783 3232
rect 4463 2144 4471 2208
rect 4535 2144 4551 2208
rect 4615 2144 4631 2208
rect 4695 2144 4711 2208
rect 4775 2144 4783 2208
rect 4463 1120 4783 2144
rect 4463 1056 4471 1120
rect 4535 1056 4551 1120
rect 4615 1056 4631 1120
rect 4695 1056 4711 1120
rect 4775 1056 4783 1120
rect 4463 496 4783 1056
rect 5820 9280 6140 9296
rect 5820 9216 5828 9280
rect 5892 9216 5908 9280
rect 5972 9216 5988 9280
rect 6052 9216 6068 9280
rect 6132 9216 6140 9280
rect 5820 8192 6140 9216
rect 5820 8128 5828 8192
rect 5892 8128 5908 8192
rect 5972 8128 5988 8192
rect 6052 8128 6068 8192
rect 6132 8128 6140 8192
rect 5820 7104 6140 8128
rect 5820 7040 5828 7104
rect 5892 7040 5908 7104
rect 5972 7040 5988 7104
rect 6052 7040 6068 7104
rect 6132 7040 6140 7104
rect 5820 6016 6140 7040
rect 5820 5952 5828 6016
rect 5892 5952 5908 6016
rect 5972 5952 5988 6016
rect 6052 5952 6068 6016
rect 6132 5952 6140 6016
rect 5820 4928 6140 5952
rect 5820 4864 5828 4928
rect 5892 4864 5908 4928
rect 5972 4864 5988 4928
rect 6052 4864 6068 4928
rect 6132 4864 6140 4928
rect 5820 3840 6140 4864
rect 5820 3776 5828 3840
rect 5892 3776 5908 3840
rect 5972 3776 5988 3840
rect 6052 3776 6068 3840
rect 6132 3776 6140 3840
rect 5820 2752 6140 3776
rect 5820 2688 5828 2752
rect 5892 2688 5908 2752
rect 5972 2688 5988 2752
rect 6052 2688 6068 2752
rect 6132 2688 6140 2752
rect 5820 1664 6140 2688
rect 5820 1600 5828 1664
rect 5892 1600 5908 1664
rect 5972 1600 5988 1664
rect 6052 1600 6068 1664
rect 6132 1600 6140 1664
rect 5820 576 6140 1600
rect 5820 512 5828 576
rect 5892 512 5908 576
rect 5972 512 5988 576
rect 6052 512 6068 576
rect 6132 512 6140 576
rect 5820 496 6140 512
rect 7177 8736 7497 9296
rect 7177 8672 7185 8736
rect 7249 8672 7265 8736
rect 7329 8672 7345 8736
rect 7409 8672 7425 8736
rect 7489 8672 7497 8736
rect 7177 7648 7497 8672
rect 7177 7584 7185 7648
rect 7249 7584 7265 7648
rect 7329 7584 7345 7648
rect 7409 7584 7425 7648
rect 7489 7584 7497 7648
rect 7177 6560 7497 7584
rect 7177 6496 7185 6560
rect 7249 6496 7265 6560
rect 7329 6496 7345 6560
rect 7409 6496 7425 6560
rect 7489 6496 7497 6560
rect 7177 5472 7497 6496
rect 8534 9280 8854 9296
rect 8534 9216 8542 9280
rect 8606 9216 8622 9280
rect 8686 9216 8702 9280
rect 8766 9216 8782 9280
rect 8846 9216 8854 9280
rect 8534 8192 8854 9216
rect 8534 8128 8542 8192
rect 8606 8128 8622 8192
rect 8686 8128 8702 8192
rect 8766 8128 8782 8192
rect 8846 8128 8854 8192
rect 8534 7104 8854 8128
rect 8534 7040 8542 7104
rect 8606 7040 8622 7104
rect 8686 7040 8702 7104
rect 8766 7040 8782 7104
rect 8846 7040 8854 7104
rect 7603 6084 7669 6085
rect 7603 6020 7604 6084
rect 7668 6020 7669 6084
rect 7603 6019 7669 6020
rect 7177 5408 7185 5472
rect 7249 5408 7265 5472
rect 7329 5408 7345 5472
rect 7409 5408 7425 5472
rect 7489 5408 7497 5472
rect 7177 4384 7497 5408
rect 7177 4320 7185 4384
rect 7249 4320 7265 4384
rect 7329 4320 7345 4384
rect 7409 4320 7425 4384
rect 7489 4320 7497 4384
rect 7177 3296 7497 4320
rect 7177 3232 7185 3296
rect 7249 3232 7265 3296
rect 7329 3232 7345 3296
rect 7409 3232 7425 3296
rect 7489 3232 7497 3296
rect 7177 2208 7497 3232
rect 7606 2549 7666 6019
rect 8534 6016 8854 7040
rect 8534 5952 8542 6016
rect 8606 5952 8622 6016
rect 8686 5952 8702 6016
rect 8766 5952 8782 6016
rect 8846 5952 8854 6016
rect 8534 4928 8854 5952
rect 8534 4864 8542 4928
rect 8606 4864 8622 4928
rect 8686 4864 8702 4928
rect 8766 4864 8782 4928
rect 8846 4864 8854 4928
rect 8534 3840 8854 4864
rect 8534 3776 8542 3840
rect 8606 3776 8622 3840
rect 8686 3776 8702 3840
rect 8766 3776 8782 3840
rect 8846 3776 8854 3840
rect 8534 2752 8854 3776
rect 8534 2688 8542 2752
rect 8606 2688 8622 2752
rect 8686 2688 8702 2752
rect 8766 2688 8782 2752
rect 8846 2688 8854 2752
rect 7603 2548 7669 2549
rect 7603 2484 7604 2548
rect 7668 2484 7669 2548
rect 7603 2483 7669 2484
rect 7177 2144 7185 2208
rect 7249 2144 7265 2208
rect 7329 2144 7345 2208
rect 7409 2144 7425 2208
rect 7489 2144 7497 2208
rect 7177 1120 7497 2144
rect 7177 1056 7185 1120
rect 7249 1056 7265 1120
rect 7329 1056 7345 1120
rect 7409 1056 7425 1120
rect 7489 1056 7497 1120
rect 7177 496 7497 1056
rect 8534 1664 8854 2688
rect 8534 1600 8542 1664
rect 8606 1600 8622 1664
rect 8686 1600 8702 1664
rect 8766 1600 8782 1664
rect 8846 1600 8854 1664
rect 8534 576 8854 1600
rect 8534 512 8542 576
rect 8606 512 8622 576
rect 8686 512 8702 576
rect 8766 512 8782 576
rect 8846 512 8854 576
rect 8534 496 8854 512
rect 9891 8736 10211 9296
rect 9891 8672 9899 8736
rect 9963 8672 9979 8736
rect 10043 8672 10059 8736
rect 10123 8672 10139 8736
rect 10203 8672 10211 8736
rect 9891 7648 10211 8672
rect 9891 7584 9899 7648
rect 9963 7584 9979 7648
rect 10043 7584 10059 7648
rect 10123 7584 10139 7648
rect 10203 7584 10211 7648
rect 9891 6560 10211 7584
rect 9891 6496 9899 6560
rect 9963 6496 9979 6560
rect 10043 6496 10059 6560
rect 10123 6496 10139 6560
rect 10203 6496 10211 6560
rect 9891 5472 10211 6496
rect 9891 5408 9899 5472
rect 9963 5408 9979 5472
rect 10043 5408 10059 5472
rect 10123 5408 10139 5472
rect 10203 5408 10211 5472
rect 9891 4384 10211 5408
rect 9891 4320 9899 4384
rect 9963 4320 9979 4384
rect 10043 4320 10059 4384
rect 10123 4320 10139 4384
rect 10203 4320 10211 4384
rect 9891 3296 10211 4320
rect 9891 3232 9899 3296
rect 9963 3232 9979 3296
rect 10043 3232 10059 3296
rect 10123 3232 10139 3296
rect 10203 3232 10211 3296
rect 9891 2208 10211 3232
rect 9891 2144 9899 2208
rect 9963 2144 9979 2208
rect 10043 2144 10059 2208
rect 10123 2144 10139 2208
rect 10203 2144 10211 2208
rect 9891 1120 10211 2144
rect 9891 1056 9899 1120
rect 9963 1056 9979 1120
rect 10043 1056 10059 1120
rect 10123 1056 10139 1120
rect 10203 1056 10211 1120
rect 9891 496 10211 1056
rect 11248 9280 11568 9296
rect 11248 9216 11256 9280
rect 11320 9216 11336 9280
rect 11400 9216 11416 9280
rect 11480 9216 11496 9280
rect 11560 9216 11568 9280
rect 11248 8192 11568 9216
rect 11248 8128 11256 8192
rect 11320 8128 11336 8192
rect 11400 8128 11416 8192
rect 11480 8128 11496 8192
rect 11560 8128 11568 8192
rect 11248 7104 11568 8128
rect 11248 7040 11256 7104
rect 11320 7040 11336 7104
rect 11400 7040 11416 7104
rect 11480 7040 11496 7104
rect 11560 7040 11568 7104
rect 11248 6016 11568 7040
rect 11248 5952 11256 6016
rect 11320 5952 11336 6016
rect 11400 5952 11416 6016
rect 11480 5952 11496 6016
rect 11560 5952 11568 6016
rect 11248 4928 11568 5952
rect 11248 4864 11256 4928
rect 11320 4864 11336 4928
rect 11400 4864 11416 4928
rect 11480 4864 11496 4928
rect 11560 4864 11568 4928
rect 11248 3840 11568 4864
rect 11248 3776 11256 3840
rect 11320 3776 11336 3840
rect 11400 3776 11416 3840
rect 11480 3776 11496 3840
rect 11560 3776 11568 3840
rect 11248 2752 11568 3776
rect 11248 2688 11256 2752
rect 11320 2688 11336 2752
rect 11400 2688 11416 2752
rect 11480 2688 11496 2752
rect 11560 2688 11568 2752
rect 11248 1664 11568 2688
rect 11248 1600 11256 1664
rect 11320 1600 11336 1664
rect 11400 1600 11416 1664
rect 11480 1600 11496 1664
rect 11560 1600 11568 1664
rect 11248 576 11568 1600
rect 11248 512 11256 576
rect 11320 512 11336 576
rect 11400 512 11416 576
rect 11480 512 11496 576
rect 11560 512 11568 576
rect 11248 496 11568 512
use sky130_fd_sc_hd__buf_2  _080_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1704896540
transform -1 0 10396 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _082_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9476 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _083_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8004 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _084_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8556 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _085_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9660 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9568 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _087_
timestamp 1704896540
transform -1 0 10580 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10488 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8372 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _090_
timestamp 1704896540
transform 1 0 7728 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8096 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8924 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _093_
timestamp 1704896540
transform -1 0 8464 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _094_
timestamp 1704896540
transform -1 0 9936 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _095_
timestamp 1704896540
transform -1 0 9936 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9108 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _097_
timestamp 1704896540
transform -1 0 8740 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _098_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9568 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _099_
timestamp 1704896540
transform -1 0 6716 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _100_
timestamp 1704896540
transform 1 0 4876 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _101_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _102_
timestamp 1704896540
transform -1 0 8188 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 1704896540
transform 1 0 8188 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp 1704896540
transform -1 0 4692 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6164 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _106_
timestamp 1704896540
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _107_
timestamp 1704896540
transform 1 0 8464 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _108_
timestamp 1704896540
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _109_
timestamp 1704896540
transform 1 0 7084 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7084 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6532 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _112_
timestamp 1704896540
transform -1 0 6532 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113_
timestamp 1704896540
transform 1 0 6808 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _114_
timestamp 1704896540
transform 1 0 7084 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 1704896540
transform 1 0 8188 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10304 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _117_
timestamp 1704896540
transform 1 0 8464 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__a22oi_1  _118_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8188 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _119_
timestamp 1704896540
transform 1 0 2300 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _120_
timestamp 1704896540
transform -1 0 4416 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _121_
timestamp 1704896540
transform 1 0 4324 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 1704896540
transform 1 0 4692 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _123_
timestamp 1704896540
transform 1 0 9108 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _124_
timestamp 1704896540
transform -1 0 9108 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _125_
timestamp 1704896540
transform -1 0 7544 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _126_
timestamp 1704896540
transform 1 0 5888 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _127_
timestamp 1704896540
transform 1 0 6532 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _128_
timestamp 1704896540
transform 1 0 5152 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _129_
timestamp 1704896540
transform 1 0 8372 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _130_
timestamp 1704896540
transform 1 0 7544 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _131_
timestamp 1704896540
transform -1 0 4232 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _132_
timestamp 1704896540
transform -1 0 3128 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _133_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2852 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _134_
timestamp 1704896540
transform 1 0 3128 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _135_
timestamp 1704896540
transform 1 0 3588 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__nor3b_4  _136_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8188 0 1 8160
box -38 -48 1418 592
use sky130_fd_sc_hd__and2b_1  _137_
timestamp 1704896540
transform 1 0 8556 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _138_
timestamp 1704896540
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _139_
timestamp 1704896540
transform 1 0 5152 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _140_
timestamp 1704896540
transform 1 0 2668 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _141_
timestamp 1704896540
transform 1 0 2944 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _142_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _143_
timestamp 1704896540
transform -1 0 1564 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _144_
timestamp 1704896540
transform 1 0 3496 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _145_
timestamp 1704896540
transform -1 0 1288 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _146_
timestamp 1704896540
transform -1 0 2300 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3128 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1704896540
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _149_
timestamp 1704896540
transform 1 0 3220 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _150_
timestamp 1704896540
transform 1 0 2300 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _151_
timestamp 1704896540
transform -1 0 4692 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _152_
timestamp 1704896540
transform -1 0 4140 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1704896540
transform -1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5428 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _155_
timestamp 1704896540
transform -1 0 4508 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1704896540
transform 1 0 3956 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _157_
timestamp 1704896540
transform -1 0 6256 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _158_
timestamp 1704896540
transform 1 0 5428 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _159_
timestamp 1704896540
transform -1 0 7268 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _160_
timestamp 1704896540
transform 1 0 5428 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _162_
timestamp 1704896540
transform 1 0 9016 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _163_
timestamp 1704896540
transform 1 0 5336 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _164_
timestamp 1704896540
transform 1 0 9200 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfbbn_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4692 0 1 4896
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _166_
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 2430 592
use sky130_fd_sc_hd__dfxtp_1  _167_
timestamp 1704896540
transform 1 0 2300 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _168_
timestamp 1704896540
transform -1 0 3128 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _169_
timestamp 1704896540
transform 1 0 1288 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _170_
timestamp 1704896540
transform 1 0 1012 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _171_
timestamp 1704896540
transform 1 0 1656 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _172_
timestamp 1704896540
transform 1 0 3312 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _173_
timestamp 1704896540
transform 1 0 3496 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _174_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4600 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _175_
timestamp 1704896540
transform 1 0 5060 0 1 1632
box -38 -48 1970 592
use sky130_fd_sc_hd__dfbbn_2  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8556 0 1 5984
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_2  _177_
timestamp 1704896540
transform 1 0 5888 0 -1 1632
box -38 -48 1970 592
use sky130_fd_sc_hd__dfbbn_1  _178_
timestamp 1704896540
transform 1 0 8464 0 1 4896
box -38 -48 2430 592
use sky130_fd_sc_hd__buf_2  _179_
timestamp 1704896540
transform 1 0 10488 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7636 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1704896540
transform -1 0 5152 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1704896540
transform 1 0 7176 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1472 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2576 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_36
timestamp 1704896540
transform 1 0 3864 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4968 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_62
timestamp 1704896540
transform 1 0 6256 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_74
timestamp 1704896540
transform 1 0 7360 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_82
timestamp 1704896540
transform 1 0 8096 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_88
timestamp 1704896540
transform 1 0 8648 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_100
timestamp 1704896540
transform 1 0 9752 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1704896540
transform 1 0 10948 0 1 544
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_15
timestamp 1704896540
transform 1 0 1932 0 -1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_40
timestamp 1704896540
transform 1 0 4232 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_52
timestamp 1704896540
transform 1 0 5336 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_86
timestamp 1704896540
transform 1 0 8464 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_98
timestamp 1704896540
transform 1 0 9568 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_102
timestamp 1704896540
transform 1 0 9936 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_107
timestamp 1704896540
transform 1 0 10396 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 1704896540
transform 1 0 10948 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_15
timestamp 1704896540
transform 1 0 1932 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2852 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3220 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_39
timestamp 1704896540
transform 1 0 4140 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_47
timestamp 1704896540
transform 1 0 4876 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_73
timestamp 1704896540
transform 1 0 7268 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 1704896540
transform 1 0 8004 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_91
timestamp 1704896540
transform 1 0 8924 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_103
timestamp 1704896540
transform 1 0 10028 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4140 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1704896540
transform 1 0 5520 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1704896540
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_62
timestamp 1704896540
transform 1 0 6256 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_74
timestamp 1704896540
transform 1 0 7360 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_86
timestamp 1704896540
transform 1 0 8464 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_98
timestamp 1704896540
transform 1 0 9568 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 1704896540
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_113
timestamp 1704896540
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_15
timestamp 1704896540
transform 1 0 1932 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1704896540
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_37
timestamp 1704896540
transform 1 0 3956 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_43
timestamp 1704896540
transform 1 0 4508 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1704896540
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_77
timestamp 1704896540
transform 1 0 7636 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_109
timestamp 1704896540
transform 1 0 10580 0 1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_15
timestamp 1704896540
transform 1 0 1932 0 -1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_35
timestamp 1704896540
transform 1 0 3772 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_47
timestamp 1704896540
transform 1 0 4876 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_67
timestamp 1704896540
transform 1 0 6716 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_75
timestamp 1704896540
transform 1 0 7452 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_81
timestamp 1704896540
transform 1 0 8004 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_99
timestamp 1704896540
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_108
timestamp 1704896540
transform 1 0 10488 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 1704896540
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_3
timestamp 1704896540
transform 1 0 828 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_11
timestamp 1704896540
transform 1 0 1564 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4324 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_48
timestamp 1704896540
transform 1 0 4968 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_56
timestamp 1704896540
transform 1 0 5704 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_61
timestamp 1704896540
transform 1 0 6164 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_69
timestamp 1704896540
transform 1 0 6900 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_89
timestamp 1704896540
transform 1 0 8740 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_102
timestamp 1704896540
transform 1 0 9936 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_114
timestamp 1704896540
transform 1 0 11040 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1704896540
transform 1 0 5796 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_61
timestamp 1704896540
transform 1 0 6164 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_65
timestamp 1704896540
transform 1 0 6532 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_71
timestamp 1704896540
transform 1 0 7084 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_83
timestamp 1704896540
transform 1 0 8188 0 -1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_95
timestamp 1704896540
transform 1 0 9292 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_107
timestamp 1704896540
transform 1 0 10396 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1704896540
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_33
timestamp 1704896540
transform 1 0 3588 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_37
timestamp 1704896540
transform 1 0 3956 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_43
timestamp 1704896540
transform 1 0 4508 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_112
timestamp 1704896540
transform 1 0 10856 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_3
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_17
timestamp 1704896540
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_30
timestamp 1704896540
transform 1 0 3312 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_57
timestamp 1704896540
transform 1 0 5796 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_68
timestamp 1704896540
transform 1 0 6808 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_86
timestamp 1704896540
transform 1 0 8464 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_94
timestamp 1704896540
transform 1 0 9200 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_100
timestamp 1704896540
transform 1 0 9752 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1704896540
transform 1 0 10948 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_56
timestamp 1704896540
transform 1 0 5704 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1704896540
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_3
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_25
timestamp 1704896540
transform 1 0 2852 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_33
timestamp 1704896540
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_40
timestamp 1704896540
transform 1 0 4232 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_44
timestamp 1704896540
transform 1 0 4600 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_86
timestamp 1704896540
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_98
timestamp 1704896540
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_102
timestamp 1704896540
transform 1 0 9936 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_108
timestamp 1704896540
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1704896540
transform 1 0 10948 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_3
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_11
timestamp 1704896540
transform 1 0 1564 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_45
timestamp 1704896540
transform 1 0 4692 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_62
timestamp 1704896540
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_72
timestamp 1704896540
transform 1 0 7176 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_99
timestamp 1704896540
transform 1 0 9660 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_111
timestamp 1704896540
transform 1 0 10764 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_45
timestamp 1704896540
transform 1 0 4692 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_49
timestamp 1704896540
transform 1 0 5060 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1704896540
transform 1 0 5796 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_92
timestamp 1704896540
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1704896540
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1704896540
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_46
timestamp 1704896540
transform 1 0 4784 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1704896540
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_91
timestamp 1704896540
transform 1 0 8924 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_112
timestamp 1704896540
transform 1 0 10856 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1704896540
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_27
timestamp 1704896540
transform 1 0 3036 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_29
timestamp 1704896540
transform 1 0 3220 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_41
timestamp 1704896540
transform 1 0 4324 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1704896540
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1704896540
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_81
timestamp 1704896540
transform 1 0 8004 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_85
timestamp 1704896540
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_97
timestamp 1704896540
transform 1 0 9476 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1704896540
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1704896540
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6440 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 3956 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform -1 0 3956 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform -1 0 3496 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform 1 0 2300 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 2300 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform -1 0 10764 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1704896540
transform -1 0 1472 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1704896540
transform 1 0 3588 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6256 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform 1 0 8372 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1704896540
transform 1 0 10856 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_16
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 11408 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_17
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 11408 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_18
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 11408 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_19
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 11408 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_20
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 11408 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_21
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 11408 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_22
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 11408 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_23
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 11408 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_24
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 11408 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_25
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 11408 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_26
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 11408 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_27
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 11408 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_28
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 11408 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_29
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 11408 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_30
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 11408 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_31
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 11408 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_33
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_34
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_35
timestamp 1704896540
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_36
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_37
timestamp 1704896540
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_38
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_39
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_40
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_41
timestamp 1704896540
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_42
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_43
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_44
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_45
timestamp 1704896540
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_46
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_47
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_48
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_49
timestamp 1704896540
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_50
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_51
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_52
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_53
timestamp 1704896540
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_54
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_55
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_56
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_57
timestamp 1704896540
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_58
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_59
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_60
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_61
timestamp 1704896540
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_62
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_63
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_64
timestamp 1704896540
transform 1 0 3128 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_65
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_66
timestamp 1704896540
transform 1 0 8280 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_67
timestamp 1704896540
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
<< labels >>
rlabel metal2 s 6060 9248 6060 9248 4 VGND
rlabel metal1 s 5980 8704 5980 8704 4 VPWR
rlabel metal1 s 5796 4046 5796 4046 4 _000_
rlabel metal1 s 8280 7514 8280 7514 4 _001_
rlabel metal1 s 5428 7990 5428 7990 4 _002_
rlabel metal1 s 9200 7514 9200 7514 4 _003_
rlabel metal2 s 6854 4828 6854 4828 4 _004_
rlabel metal2 s 8234 6188 8234 6188 4 _005_
rlabel metal2 s 10258 4284 10258 4284 4 _006_
rlabel metal1 s 6854 5134 6854 5134 4 _007_
rlabel metal1 s 6256 4794 6256 4794 4 _008_
rlabel metal2 s 4278 5984 4278 5984 4 _009_
rlabel metal2 s 7682 6630 7682 6630 4 _010_
rlabel metal1 s 7689 6902 7689 6902 4 _011_
rlabel metal2 s 5290 6596 5290 6596 4 _012_
rlabel metal1 s 6118 3910 6118 3910 4 _013_
rlabel metal1 s 6164 2278 6164 2278 4 _014_
rlabel metal1 s 9752 6630 9752 6630 4 _015_
rlabel metal1 s 7774 6120 7774 6120 4 _016_
rlabel metal1 s 7176 1734 7176 1734 4 _017_
rlabel metal2 s 9614 5304 9614 5304 4 _018_
rlabel metal2 s 8510 5372 8510 5372 4 _019_
rlabel metal1 s 4830 5270 4830 5270 4 _020_
rlabel metal2 s 6578 6324 6578 6324 4 _021_
rlabel metal1 s 2668 3162 2668 3162 4 _022_
rlabel metal1 s 2810 4046 2810 4046 4 _023_
rlabel metal1 s 1242 4794 1242 4794 4 _024_
rlabel metal2 s 1329 6222 1329 6222 4 _025_
rlabel metal2 s 2346 7106 2346 7106 4 _026_
rlabel metal1 s 3542 7786 3542 7786 4 _027_
rlabel metal1 s 3905 5814 3905 5814 4 _028_
rlabel metal2 s 4922 3196 4922 3196 4 _029_
rlabel metal2 s 5382 2108 5382 2108 4 _030_
rlabel metal1 s 9246 4114 9246 4114 4 _031_
rlabel metal1 s 7866 1292 7866 1292 4 _032_
rlabel metal2 s 8418 4386 8418 4386 4 _033_
rlabel metal2 s 9706 3876 9706 3876 4 _034_
rlabel metal1 s 8326 4794 8326 4794 4 _035_
rlabel metal1 s 3772 6834 3772 6834 4 _036_
rlabel metal1 s 4048 7514 4048 7514 4 _037_
rlabel metal1 s 8418 7276 8418 7276 4 _038_
rlabel metal2 s 6394 7616 6394 7616 4 _039_
rlabel metal1 s 5796 7854 5796 7854 4 _040_
rlabel metal2 s 6578 7650 6578 7650 4 _041_
rlabel metal1 s 8280 7310 8280 7310 4 _042_
rlabel metal1 s 3634 1496 3634 1496 4 _043_
rlabel metal2 s 2714 1666 2714 1666 4 _044_
rlabel metal2 s 3542 1666 3542 1666 4 _045_
rlabel metal1 s 9154 8976 9154 8976 4 _046_
rlabel metal1 s 3220 5134 3220 5134 4 _047_
rlabel metal1 s 2162 5236 2162 5236 4 _048_
rlabel metal1 s 2392 4658 2392 4658 4 _049_
rlabel metal1 s 2484 6426 2484 6426 4 _050_
rlabel metal1 s 2530 6324 2530 6324 4 _051_
rlabel metal1 s 2530 6766 2530 6766 4 _052_
rlabel metal1 s 4186 7718 4186 7718 4 _053_
rlabel metal1 s 3404 7922 3404 7922 4 _054_
rlabel metal1 s 4638 4998 4638 4998 4 _055_
rlabel metal1 s 4140 5338 4140 5338 4 _056_
rlabel metal1 s 4600 5066 4600 5066 4 _057_
rlabel metal1 s 6256 4046 6256 4046 4 _058_
rlabel metal1 s 8694 3502 8694 3502 4 _059_
rlabel metal1 s 9246 2992 9246 2992 4 _060_
rlabel metal1 s 6670 3434 6670 3434 4 _061_
rlabel metal2 s 8878 4012 8878 4012 4 _062_
rlabel metal2 s 10442 3332 10442 3332 4 _063_
rlabel metal1 s 9062 3434 9062 3434 4 _064_
rlabel metal2 s 7774 3366 7774 3366 4 _065_
rlabel metal1 s 6394 3434 6394 3434 4 _066_
rlabel metal1 s 8280 1326 8280 1326 4 _067_
rlabel metal2 s 9154 4352 9154 4352 4 _068_
rlabel metal1 s 9108 3706 9108 3706 4 _069_
rlabel metal1 s 8878 4012 8878 4012 4 _070_
rlabel metal1 s 5888 3570 5888 3570 4 _071_
rlabel metal2 s 8326 6052 8326 6052 4 _072_
rlabel metal1 s 8326 3706 8326 3706 4 _073_
rlabel metal1 s 7958 5168 7958 5168 4 _074_
rlabel metal2 s 7771 5134 7771 5134 4 _075_
rlabel metal1 s 6831 5746 6831 5746 4 _076_
rlabel metal1 s 7222 4794 7222 4794 4 _077_
rlabel metal1 s 8372 6630 8372 6630 4 _078_
rlabel metal2 s 1150 568 1150 568 4 analog_to_digital_in[0]
rlabel metal2 s 3542 568 3542 568 4 analog_to_digital_in[1]
rlabel metal2 s 5906 0 5962 400 4 analog_to_digital_in[2]
port 5 nsew
rlabel metal2 s 8326 568 8326 568 4 analog_to_digital_in[3]
rlabel metal2 s 10718 874 10718 874 4 btn
rlabel metal2 s 7590 6103 7590 6103 4 clk
rlabel metal1 s 6578 6426 6578 6426 4 clknet_0_clk
rlabel metal1 s 3036 4046 3036 4046 4 clknet_1_0__leaf_clk
rlabel metal1 s 5106 8398 5106 8398 4 clknet_1_1__leaf_clk
rlabel metal1 s 6762 8330 6762 8330 4 control[0]
rlabel metal1 s 8832 9146 8832 9146 4 control[1]
rlabel metal2 s 10718 9156 10718 9156 4 control[2]
rlabel metal1 s 1978 2074 1978 2074 4 encoded_out[0]
rlabel metal2 s 3641 9724 3641 9724 4 encoded_out[1]
rlabel metal2 s 1426 1190 1426 1190 4 net1
rlabel metal1 s 2254 5066 2254 5066 4 net10
rlabel metal1 s 1058 4692 1058 4692 4 net11
rlabel metal2 s 1605 4726 1605 4726 4 net12
rlabel metal1 s 9338 7276 9338 7276 4 net13
rlabel metal2 s 3358 1088 3358 1088 4 net2
rlabel metal1 s 4784 1394 4784 1394 4 net3
rlabel metal2 s 4094 1122 4094 1122 4 net4
rlabel metal2 s 10442 5678 10442 5678 4 net5
rlabel metal2 s 7038 7548 7038 7548 4 net6
rlabel metal1 s 3496 5134 3496 5134 4 net7
rlabel metal1 s 3542 6970 3542 6970 4 net8
rlabel metal2 s 2806 4964 2806 4964 4 net9
rlabel metal2 s 11086 7361 11086 7361 4 reset_n
rlabel metal1 s 6348 7514 6348 7514 4 traffic_lights.control_unit.state_traffic_lights\[0\]
rlabel metal2 s 8970 8738 8970 8738 4 traffic_lights.control_unit.state_traffic_lights\[1\]
rlabel metal2 s 6762 8092 6762 8092 4 traffic_lights.control_unit.state_traffic_lights\[2\]
rlabel metal1 s 6762 7242 6762 7242 4 traffic_lights.control_unit.state_traffic_lights\[3\]
rlabel metal1 s 6302 4692 6302 4692 4 traffic_lights.control_unit.sw_traffic_lights\[0\]
rlabel metal1 s 7682 5882 7682 5882 4 traffic_lights.control_unit.sw_traffic_lights\[1\]
rlabel metal1 s 2668 5882 2668 5882 4 traffic_lights.datapath.counter.processQ\[0\]
rlabel metal1 s 2162 5746 2162 5746 4 traffic_lights.datapath.counter.processQ\[1\]
rlabel metal1 s 2346 5882 2346 5882 4 traffic_lights.datapath.counter.processQ\[2\]
rlabel metal1 s 2300 6358 2300 6358 4 traffic_lights.datapath.counter.processQ\[3\]
rlabel metal1 s 3818 7412 3818 7412 4 traffic_lights.datapath.counter.processQ\[4\]
rlabel metal1 s 4600 7922 4600 7922 4 traffic_lights.datapath.counter.processQ\[5\]
rlabel metal2 s 4922 6358 4922 6358 4 traffic_lights.datapath.counter.processQ\[6\]
rlabel metal1 s 4646 2924 4646 2924 4 traffic_lights.datapath.counter.roll
rlabel metal1 s 6394 2992 6394 2992 4 traffic_lights.datapath.glue_logic.time_length\[0\]
rlabel metal1 s 8924 3026 8924 3026 4 traffic_lights.datapath.glue_logic.time_length\[1\]
rlabel metal2 s 9798 5168 9798 5168 4 traffic_lights.datapath.glue_logic.time_length\[2\]
rlabel metal2 s 8878 3026 8878 3026 4 traffic_lights.datapath.glue_logic.time_length\[3\]
rlabel metal2 s 9614 4131 9614 4131 4 traffic_lights.datapath.glue_logic.time_length\[4\]
flabel metal4 s 11248 496 11568 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 8534 496 8854 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5820 496 6140 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3106 496 3426 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 9891 496 10211 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7177 496 7497 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4463 496 4783 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1749 496 2069 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 1122 0 1178 400 0 FreeSans 280 90 0 0 analog_to_digital_in[0]
port 3 nsew
flabel metal2 s 3514 0 3570 400 0 FreeSans 280 90 0 0 analog_to_digital_in[1]
port 4 nsew
flabel metal2 s 5934 200 5934 200 0 FreeSans 280 90 0 0 analog_to_digital_in[2]
flabel metal2 s 8298 0 8354 400 0 FreeSans 280 90 0 0 analog_to_digital_in[3]
port 6 nsew
flabel metal2 s 10690 0 10746 400 0 FreeSans 280 90 0 0 btn
port 7 nsew
flabel metal3 s 11600 2456 12000 2576 0 FreeSans 600 0 0 0 clk
port 8 nsew
flabel metal2 s 5906 9600 5962 10000 0 FreeSans 280 90 0 0 control[0]
port 9 nsew
flabel metal2 s 8298 9600 8354 10000 0 FreeSans 280 90 0 0 control[1]
port 10 nsew
flabel metal2 s 10690 9600 10746 10000 0 FreeSans 280 90 0 0 control[2]
port 11 nsew
flabel metal2 s 1122 9600 1178 10000 0 FreeSans 280 90 0 0 encoded_out[0]
port 12 nsew
flabel metal2 s 3514 9600 3570 10000 0 FreeSans 280 90 0 0 encoded_out[1]
port 13 nsew
flabel metal3 s 11600 7352 12000 7472 0 FreeSans 600 0 0 0 reset_n
port 14 nsew
<< properties >>
string FIXED_BBOX 0 0 12000 10000
string GDS_END 551996
string GDS_FILE ../gds/adc_digital_control.gds
string GDS_START 239470
<< end >>
