magic
tech sky130A
magscale 1 2
timestamp 1728848001
<< viali >>
rect -416 2304 -382 2510
rect -588 2216 -382 2250
rect -1672 760 110 794
<< metal1 >>
rect 2328 6013 2528 6050
rect 2328 5883 2362 6013
rect 2492 5883 2528 6013
rect 2328 5850 2528 5883
rect 4818 6013 5018 6050
rect 4818 5883 4854 6013
rect 4984 5883 5018 6013
rect 4818 5850 5018 5883
rect 7310 6019 7510 6050
rect 7310 5889 7346 6019
rect 7476 5889 7510 6019
rect 7310 5850 7510 5889
rect 9804 6017 10004 6050
rect 9804 5887 9838 6017
rect 9968 5887 10004 6017
rect 9804 5850 10004 5887
rect -1708 5450 806 5650
rect -286 4302 -148 5450
rect 2362 5303 2492 5309
rect 2362 3823 2492 5173
rect 4854 5303 4984 5309
rect 4854 3501 4984 5173
rect 7346 5303 7476 5309
rect 7346 3763 7476 5173
rect 9838 5303 9968 5309
rect 9838 4177 9968 5173
rect -1534 2486 -1334 2544
rect -1534 2398 -1476 2486
rect -1388 2398 -1334 2486
rect -1534 2344 -1334 2398
rect -422 2510 -370 2522
rect -422 2304 -416 2510
rect -382 2304 -370 2510
rect -422 2256 -370 2304
rect -600 2250 -370 2256
rect -600 2216 -588 2250
rect -382 2216 -370 2250
rect -600 2210 -370 2216
rect -286 2272 -148 2866
rect -286 2184 -260 2272
rect -172 2184 -148 2272
rect -286 2120 -148 2184
rect 252 2272 340 2278
rect 252 2178 340 2184
rect 2744 2272 2832 2278
rect 2744 2178 2832 2184
rect 5237 2272 5327 2278
rect 5237 2176 5327 2182
rect 7728 2270 7816 2276
rect 7728 2176 7816 2182
rect -1542 1938 -1110 2120
rect -452 1982 -20 2120
rect -1542 1800 -20 1938
rect -1542 1576 -1110 1756
rect -452 1732 -20 1800
rect -452 1644 -144 1732
rect -56 1644 -20 1732
rect -452 1618 -20 1644
rect -1542 1438 -20 1576
rect -1542 1212 -1110 1392
rect -452 1366 -20 1438
rect -452 1278 -144 1366
rect -56 1278 -20 1366
rect -452 1254 -20 1278
rect -1542 1074 -20 1212
rect -1542 800 -1110 1028
rect -452 1004 -20 1074
rect -452 916 -144 1004
rect -56 916 -20 1004
rect -452 890 -20 916
rect -1708 794 200 800
rect -1708 760 -1672 794
rect 110 760 200 794
rect -1708 600 200 760
rect 202 600 402 800
rect 488 600 630 800
<< via1 >>
rect 2362 5883 2492 6013
rect 4854 5883 4984 6013
rect 7346 5889 7476 6019
rect 9838 5887 9968 6017
rect 2362 5173 2492 5303
rect 4854 5173 4984 5303
rect 7346 5173 7476 5303
rect 9838 5173 9968 5303
rect -1476 2398 -1388 2486
rect -260 2184 -172 2272
rect 252 2184 340 2272
rect 2744 2184 2832 2272
rect 5237 2182 5327 2272
rect 7728 2182 7816 2270
rect -144 1644 -56 1732
rect -144 1278 -56 1366
rect -144 916 -56 1004
<< metal2 >>
rect 7346 6019 7476 6025
rect 2362 6013 2492 6019
rect 2362 5303 2492 5883
rect 4854 6013 4984 6019
rect 4854 5303 4984 5883
rect 7346 5303 7476 5889
rect 9838 6017 9968 6023
rect 9838 5303 9968 5887
rect 2356 5173 2362 5303
rect 2492 5173 2498 5303
rect 4848 5173 4854 5303
rect 4984 5173 4990 5303
rect 7340 5173 7346 5303
rect 7476 5173 7482 5303
rect 9832 5173 9838 5303
rect 9968 5173 9974 5303
rect -951 2486 -873 2490
rect -1482 2398 -1476 2486
rect -1388 2481 -868 2486
rect -1388 2403 -951 2481
rect -873 2403 -868 2481
rect -1388 2398 -868 2403
rect -951 2394 -873 2398
rect -266 2184 -260 2272
rect -172 2184 252 2272
rect 340 2184 346 2272
rect 2534 2184 2744 2272
rect 2832 2184 2838 2272
rect 5104 2270 5237 2272
rect 2534 1732 2622 2184
rect -150 1644 -144 1732
rect -56 1730 0 1732
rect 200 1730 2622 1732
rect -56 1644 2622 1730
rect 5020 2182 5237 2270
rect 5327 2182 5333 2272
rect 7514 2182 7728 2270
rect 7816 2182 7822 2270
rect 5020 1366 5108 2182
rect -150 1278 -144 1366
rect -56 1278 5108 1366
rect 7514 1004 7602 2182
rect -150 916 -144 1004
rect -56 916 7602 1004
<< via2 >>
rect -951 2403 -873 2481
<< metal3 >>
rect -956 2481 9352 2486
rect -956 2403 -951 2481
rect -873 2403 9352 2481
rect -956 2398 9352 2403
rect 440 2334 1600 2398
rect 2932 2334 4092 2398
rect 5424 2334 6584 2398
rect 7916 2334 9076 2398
use opamp  x1
timestamp 1728846299
transform 1 0 928 0 1 1928
box 6548 -1328 9040 3722
use opamp  x2
timestamp 1728846299
transform 1 0 -1564 0 1 1928
box 6548 -1328 9040 3722
use opamp  x3
timestamp 1728846299
transform 1 0 -4056 0 1 1928
box 6548 -1328 9040 3722
use opamp  x4
timestamp 1728846299
transform 1 0 -6548 0 1 1928
box 6548 -1328 9040 3722
use sky130_fd_pr__res_high_po_0p69_PFVE8M  XR1
timestamp 1728801405
transform -1 0 -217 0 -1 3584
box -235 -1316 235 1316
use sky130_fd_pr__res_high_po_0p69_B9B9MH  XR2
timestamp 1728801405
transform 0 1 -781 -1 0 2051
box -235 -927 235 927
use sky130_fd_pr__res_high_po_0p69_B9B9MH  XR3
timestamp 1728801405
transform 0 1 -781 -1 0 1687
box -235 -927 235 927
use sky130_fd_pr__res_high_po_0p69_B9B9MH  XR4
timestamp 1728801405
transform 0 1 -781 -1 0 1323
box -235 -927 235 927
use sky130_fd_pr__res_high_po_0p69_B9B9MH  XR5
timestamp 1728801405
transform 0 1 -781 -1 0 959
box -235 -927 235 927
<< labels >>
flabel metal1 202 5450 402 5650 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 202 600 402 800 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 2328 5850 2528 6050 0 FreeSans 256 0 0 0 out3
port 3 nsew
flabel metal1 4818 5850 5018 6050 0 FreeSans 256 0 0 0 out2
port 4 nsew
flabel metal1 7310 5850 7510 6050 0 FreeSans 256 0 0 0 out1
port 5 nsew
flabel metal1 9804 5850 10004 6050 0 FreeSans 256 0 0 0 out0
port 6 nsew
flabel metal1 -1534 2344 -1334 2544 0 FreeSans 256 0 0 0 in
port 1 nsew
<< end >>
