magic
tech sky130A
magscale 1 2
timestamp 1727826562
<< viali >>
rect 1987 1513 2021 1547
rect 2237 1513 2271 1547
rect 3249 1513 3283 1547
rect 3525 1513 3559 1547
rect 1777 1445 1811 1479
rect 2881 1445 2915 1479
rect 3081 1445 3115 1479
rect 2605 1377 2639 1411
rect 3341 1377 3375 1411
rect 2697 1309 2731 1343
rect 1961 1173 1995 1207
rect 2145 1173 2179 1207
rect 3065 1173 3099 1207
rect 2053 969 2087 1003
rect 2513 969 2547 1003
rect 3249 969 3283 1003
rect 1041 901 1075 935
rect 3893 901 3927 935
rect 857 765 891 799
rect 2237 765 2271 799
rect 2329 765 2363 799
rect 3433 765 3467 799
rect 4077 765 4111 799
<< metal1 >>
rect 552 2202 4416 2224
rect 552 2150 881 2202
rect 933 2150 945 2202
rect 997 2150 1009 2202
rect 1061 2150 1073 2202
rect 1125 2150 1137 2202
rect 1189 2150 1847 2202
rect 1899 2150 1911 2202
rect 1963 2150 1975 2202
rect 2027 2150 2039 2202
rect 2091 2150 2103 2202
rect 2155 2150 2813 2202
rect 2865 2150 2877 2202
rect 2929 2150 2941 2202
rect 2993 2150 3005 2202
rect 3057 2150 3069 2202
rect 3121 2150 3779 2202
rect 3831 2150 3843 2202
rect 3895 2150 3907 2202
rect 3959 2150 3971 2202
rect 4023 2150 4035 2202
rect 4087 2150 4416 2202
rect 552 2128 4416 2150
rect 552 1658 4576 1680
rect 552 1606 1364 1658
rect 1416 1606 1428 1658
rect 1480 1606 1492 1658
rect 1544 1606 1556 1658
rect 1608 1606 1620 1658
rect 1672 1606 2330 1658
rect 2382 1606 2394 1658
rect 2446 1606 2458 1658
rect 2510 1606 2522 1658
rect 2574 1606 2586 1658
rect 2638 1606 3296 1658
rect 3348 1606 3360 1658
rect 3412 1606 3424 1658
rect 3476 1606 3488 1658
rect 3540 1606 3552 1658
rect 3604 1606 4262 1658
rect 4314 1606 4326 1658
rect 4378 1606 4390 1658
rect 4442 1606 4454 1658
rect 4506 1606 4518 1658
rect 4570 1606 4576 1658
rect 552 1584 4576 1606
rect 1975 1547 2033 1553
rect 1975 1513 1987 1547
rect 2021 1544 2033 1547
rect 2225 1547 2283 1553
rect 2225 1544 2237 1547
rect 2021 1516 2237 1544
rect 2021 1513 2033 1516
rect 1975 1507 2033 1513
rect 2225 1513 2237 1516
rect 2271 1513 2283 1547
rect 2225 1507 2283 1513
rect 3237 1547 3295 1553
rect 3237 1513 3249 1547
rect 3283 1513 3295 1547
rect 3237 1507 3295 1513
rect 3513 1547 3571 1553
rect 3513 1513 3525 1547
rect 3559 1544 3571 1547
rect 3694 1544 3700 1556
rect 3559 1516 3700 1544
rect 3559 1513 3571 1516
rect 3513 1507 3571 1513
rect 1765 1479 1823 1485
rect 1765 1445 1777 1479
rect 1811 1476 1823 1479
rect 2498 1476 2504 1488
rect 1811 1448 2504 1476
rect 1811 1445 1823 1448
rect 1765 1439 1823 1445
rect 2498 1436 2504 1448
rect 2556 1476 2562 1488
rect 2869 1479 2927 1485
rect 2869 1476 2881 1479
rect 2556 1448 2881 1476
rect 2556 1436 2562 1448
rect 2869 1445 2881 1448
rect 2915 1445 2927 1479
rect 3069 1479 3127 1485
rect 3069 1476 3081 1479
rect 2869 1439 2927 1445
rect 3068 1445 3081 1476
rect 3115 1445 3127 1479
rect 3068 1439 3127 1445
rect 2590 1368 2596 1420
rect 2648 1368 2654 1420
rect 2685 1343 2743 1349
rect 2685 1309 2697 1343
rect 2731 1340 2743 1343
rect 3068 1340 3096 1439
rect 3252 1408 3280 1507
rect 3694 1504 3700 1516
rect 3752 1504 3758 1556
rect 3329 1411 3387 1417
rect 3329 1408 3341 1411
rect 3252 1380 3341 1408
rect 3329 1377 3341 1380
rect 3375 1377 3387 1411
rect 3329 1371 3387 1377
rect 3234 1340 3240 1352
rect 2731 1312 3240 1340
rect 2731 1309 2743 1312
rect 2685 1303 2743 1309
rect 3234 1300 3240 1312
rect 3292 1300 3298 1352
rect 1964 1244 3096 1272
rect 1762 1164 1768 1216
rect 1820 1204 1826 1216
rect 1964 1213 1992 1244
rect 1949 1207 2007 1213
rect 1949 1204 1961 1207
rect 1820 1176 1961 1204
rect 1820 1164 1826 1176
rect 1949 1173 1961 1176
rect 1995 1173 2007 1207
rect 1949 1167 2007 1173
rect 2133 1207 2191 1213
rect 2133 1173 2145 1207
rect 2179 1204 2191 1207
rect 2222 1204 2228 1216
rect 2179 1176 2228 1204
rect 2179 1173 2191 1176
rect 2133 1167 2191 1173
rect 2222 1164 2228 1176
rect 2280 1164 2286 1216
rect 3068 1213 3096 1244
rect 3053 1207 3111 1213
rect 3053 1173 3065 1207
rect 3099 1173 3111 1207
rect 3053 1167 3111 1173
rect 552 1114 4416 1136
rect 552 1062 881 1114
rect 933 1062 945 1114
rect 997 1062 1009 1114
rect 1061 1062 1073 1114
rect 1125 1062 1137 1114
rect 1189 1062 1847 1114
rect 1899 1062 1911 1114
rect 1963 1062 1975 1114
rect 2027 1062 2039 1114
rect 2091 1062 2103 1114
rect 2155 1062 2813 1114
rect 2865 1062 2877 1114
rect 2929 1062 2941 1114
rect 2993 1062 3005 1114
rect 3057 1062 3069 1114
rect 3121 1062 3779 1114
rect 3831 1062 3843 1114
rect 3895 1062 3907 1114
rect 3959 1062 3971 1114
rect 4023 1062 4035 1114
rect 4087 1062 4416 1114
rect 552 1040 4416 1062
rect 1210 960 1216 1012
rect 1268 1000 1274 1012
rect 2041 1003 2099 1009
rect 2041 1000 2053 1003
rect 1268 972 2053 1000
rect 1268 960 1274 972
rect 2041 969 2053 972
rect 2087 969 2099 1003
rect 2041 963 2099 969
rect 2498 960 2504 1012
rect 2556 960 2562 1012
rect 3234 960 3240 1012
rect 3292 960 3298 1012
rect 1029 935 1087 941
rect 1029 901 1041 935
rect 1075 932 1087 935
rect 1762 932 1768 944
rect 1075 904 1768 932
rect 1075 901 1087 904
rect 1029 895 1087 901
rect 1762 892 1768 904
rect 1820 892 1826 944
rect 2590 892 2596 944
rect 2648 932 2654 944
rect 3881 935 3939 941
rect 3881 932 3893 935
rect 2648 904 3893 932
rect 2648 892 2654 904
rect 3881 901 3893 904
rect 3927 901 3939 935
rect 3881 895 3939 901
rect 658 756 664 808
rect 716 796 722 808
rect 845 799 903 805
rect 845 796 857 799
rect 716 768 857 796
rect 716 756 722 768
rect 845 765 857 768
rect 891 765 903 799
rect 845 759 903 765
rect 2222 756 2228 808
rect 2280 756 2286 808
rect 2317 799 2375 805
rect 2317 765 2329 799
rect 2363 765 2375 799
rect 2317 759 2375 765
rect 1854 688 1860 740
rect 1912 728 1918 740
rect 2332 728 2360 759
rect 3050 756 3056 808
rect 3108 796 3114 808
rect 3421 799 3479 805
rect 3421 796 3433 799
rect 3108 768 3433 796
rect 3108 756 3114 768
rect 3421 765 3433 768
rect 3467 765 3479 799
rect 3421 759 3479 765
rect 4062 756 4068 808
rect 4120 756 4126 808
rect 1912 700 2360 728
rect 1912 688 1918 700
rect 552 570 4576 592
rect 552 518 1364 570
rect 1416 518 1428 570
rect 1480 518 1492 570
rect 1544 518 1556 570
rect 1608 518 1620 570
rect 1672 518 2330 570
rect 2382 518 2394 570
rect 2446 518 2458 570
rect 2510 518 2522 570
rect 2574 518 2586 570
rect 2638 518 3296 570
rect 3348 518 3360 570
rect 3412 518 3424 570
rect 3476 518 3488 570
rect 3540 518 3552 570
rect 3604 518 4262 570
rect 4314 518 4326 570
rect 4378 518 4390 570
rect 4442 518 4454 570
rect 4506 518 4518 570
rect 4570 518 4576 570
rect 552 496 4576 518
rect 4062 416 4068 468
rect 4120 456 4126 468
rect 4338 456 4344 468
rect 4120 428 4344 456
rect 4120 416 4126 428
rect 4338 416 4344 428
rect 4396 416 4402 468
<< via1 >>
rect 881 2150 933 2202
rect 945 2150 997 2202
rect 1009 2150 1061 2202
rect 1073 2150 1125 2202
rect 1137 2150 1189 2202
rect 1847 2150 1899 2202
rect 1911 2150 1963 2202
rect 1975 2150 2027 2202
rect 2039 2150 2091 2202
rect 2103 2150 2155 2202
rect 2813 2150 2865 2202
rect 2877 2150 2929 2202
rect 2941 2150 2993 2202
rect 3005 2150 3057 2202
rect 3069 2150 3121 2202
rect 3779 2150 3831 2202
rect 3843 2150 3895 2202
rect 3907 2150 3959 2202
rect 3971 2150 4023 2202
rect 4035 2150 4087 2202
rect 1364 1606 1416 1658
rect 1428 1606 1480 1658
rect 1492 1606 1544 1658
rect 1556 1606 1608 1658
rect 1620 1606 1672 1658
rect 2330 1606 2382 1658
rect 2394 1606 2446 1658
rect 2458 1606 2510 1658
rect 2522 1606 2574 1658
rect 2586 1606 2638 1658
rect 3296 1606 3348 1658
rect 3360 1606 3412 1658
rect 3424 1606 3476 1658
rect 3488 1606 3540 1658
rect 3552 1606 3604 1658
rect 4262 1606 4314 1658
rect 4326 1606 4378 1658
rect 4390 1606 4442 1658
rect 4454 1606 4506 1658
rect 4518 1606 4570 1658
rect 2504 1436 2556 1488
rect 2596 1411 2648 1420
rect 2596 1377 2605 1411
rect 2605 1377 2639 1411
rect 2639 1377 2648 1411
rect 2596 1368 2648 1377
rect 3700 1504 3752 1556
rect 3240 1300 3292 1352
rect 1768 1164 1820 1216
rect 2228 1164 2280 1216
rect 881 1062 933 1114
rect 945 1062 997 1114
rect 1009 1062 1061 1114
rect 1073 1062 1125 1114
rect 1137 1062 1189 1114
rect 1847 1062 1899 1114
rect 1911 1062 1963 1114
rect 1975 1062 2027 1114
rect 2039 1062 2091 1114
rect 2103 1062 2155 1114
rect 2813 1062 2865 1114
rect 2877 1062 2929 1114
rect 2941 1062 2993 1114
rect 3005 1062 3057 1114
rect 3069 1062 3121 1114
rect 3779 1062 3831 1114
rect 3843 1062 3895 1114
rect 3907 1062 3959 1114
rect 3971 1062 4023 1114
rect 4035 1062 4087 1114
rect 1216 960 1268 1012
rect 2504 1003 2556 1012
rect 2504 969 2513 1003
rect 2513 969 2547 1003
rect 2547 969 2556 1003
rect 2504 960 2556 969
rect 3240 1003 3292 1012
rect 3240 969 3249 1003
rect 3249 969 3283 1003
rect 3283 969 3292 1003
rect 3240 960 3292 969
rect 1768 892 1820 944
rect 2596 892 2648 944
rect 664 756 716 808
rect 2228 799 2280 808
rect 2228 765 2237 799
rect 2237 765 2271 799
rect 2271 765 2280 799
rect 2228 756 2280 765
rect 1860 688 1912 740
rect 3056 756 3108 808
rect 4068 799 4120 808
rect 4068 765 4077 799
rect 4077 765 4111 799
rect 4111 765 4120 799
rect 4068 756 4120 765
rect 1364 518 1416 570
rect 1428 518 1480 570
rect 1492 518 1544 570
rect 1556 518 1608 570
rect 1620 518 1672 570
rect 2330 518 2382 570
rect 2394 518 2446 570
rect 2458 518 2510 570
rect 2522 518 2574 570
rect 2586 518 2638 570
rect 3296 518 3348 570
rect 3360 518 3412 570
rect 3424 518 3476 570
rect 3488 518 3540 570
rect 3552 518 3604 570
rect 4262 518 4314 570
rect 4326 518 4378 570
rect 4390 518 4442 570
rect 4454 518 4506 570
rect 4518 518 4570 570
rect 4068 416 4120 468
rect 4344 416 4396 468
<< metal2 >>
rect 1214 2600 1270 3000
rect 3698 2600 3754 3000
rect 881 2204 1189 2213
rect 881 2202 887 2204
rect 943 2202 967 2204
rect 1023 2202 1047 2204
rect 1103 2202 1127 2204
rect 1183 2202 1189 2204
rect 943 2150 945 2202
rect 1125 2150 1127 2202
rect 881 2148 887 2150
rect 943 2148 967 2150
rect 1023 2148 1047 2150
rect 1103 2148 1127 2150
rect 1183 2148 1189 2150
rect 881 2139 1189 2148
rect 881 1116 1189 1125
rect 881 1114 887 1116
rect 943 1114 967 1116
rect 1023 1114 1047 1116
rect 1103 1114 1127 1116
rect 1183 1114 1189 1116
rect 943 1062 945 1114
rect 1125 1062 1127 1114
rect 881 1060 887 1062
rect 943 1060 967 1062
rect 1023 1060 1047 1062
rect 1103 1060 1127 1062
rect 1183 1060 1189 1062
rect 881 1051 1189 1060
rect 1228 1018 1256 2600
rect 1847 2204 2155 2213
rect 1847 2202 1853 2204
rect 1909 2202 1933 2204
rect 1989 2202 2013 2204
rect 2069 2202 2093 2204
rect 2149 2202 2155 2204
rect 1909 2150 1911 2202
rect 2091 2150 2093 2202
rect 1847 2148 1853 2150
rect 1909 2148 1933 2150
rect 1989 2148 2013 2150
rect 2069 2148 2093 2150
rect 2149 2148 2155 2150
rect 1847 2139 2155 2148
rect 2813 2204 3121 2213
rect 2813 2202 2819 2204
rect 2875 2202 2899 2204
rect 2955 2202 2979 2204
rect 3035 2202 3059 2204
rect 3115 2202 3121 2204
rect 2875 2150 2877 2202
rect 3057 2150 3059 2202
rect 2813 2148 2819 2150
rect 2875 2148 2899 2150
rect 2955 2148 2979 2150
rect 3035 2148 3059 2150
rect 3115 2148 3121 2150
rect 2813 2139 3121 2148
rect 1364 1660 1672 1669
rect 1364 1658 1370 1660
rect 1426 1658 1450 1660
rect 1506 1658 1530 1660
rect 1586 1658 1610 1660
rect 1666 1658 1672 1660
rect 1426 1606 1428 1658
rect 1608 1606 1610 1658
rect 1364 1604 1370 1606
rect 1426 1604 1450 1606
rect 1506 1604 1530 1606
rect 1586 1604 1610 1606
rect 1666 1604 1672 1606
rect 1364 1595 1672 1604
rect 2330 1660 2638 1669
rect 2330 1658 2336 1660
rect 2392 1658 2416 1660
rect 2472 1658 2496 1660
rect 2552 1658 2576 1660
rect 2632 1658 2638 1660
rect 2392 1606 2394 1658
rect 2574 1606 2576 1658
rect 2330 1604 2336 1606
rect 2392 1604 2416 1606
rect 2472 1604 2496 1606
rect 2552 1604 2576 1606
rect 2632 1604 2638 1606
rect 2330 1595 2638 1604
rect 3296 1660 3604 1669
rect 3296 1658 3302 1660
rect 3358 1658 3382 1660
rect 3438 1658 3462 1660
rect 3518 1658 3542 1660
rect 3598 1658 3604 1660
rect 3358 1606 3360 1658
rect 3540 1606 3542 1658
rect 3296 1604 3302 1606
rect 3358 1604 3382 1606
rect 3438 1604 3462 1606
rect 3518 1604 3542 1606
rect 3598 1604 3604 1606
rect 3296 1595 3604 1604
rect 3712 1562 3740 2600
rect 3779 2204 4087 2213
rect 3779 2202 3785 2204
rect 3841 2202 3865 2204
rect 3921 2202 3945 2204
rect 4001 2202 4025 2204
rect 4081 2202 4087 2204
rect 3841 2150 3843 2202
rect 4023 2150 4025 2202
rect 3779 2148 3785 2150
rect 3841 2148 3865 2150
rect 3921 2148 3945 2150
rect 4001 2148 4025 2150
rect 4081 2148 4087 2150
rect 3779 2139 4087 2148
rect 4262 1660 4570 1669
rect 4262 1658 4268 1660
rect 4324 1658 4348 1660
rect 4404 1658 4428 1660
rect 4484 1658 4508 1660
rect 4564 1658 4570 1660
rect 4324 1606 4326 1658
rect 4506 1606 4508 1658
rect 4262 1604 4268 1606
rect 4324 1604 4348 1606
rect 4404 1604 4428 1606
rect 4484 1604 4508 1606
rect 4564 1604 4570 1606
rect 4262 1595 4570 1604
rect 3700 1556 3752 1562
rect 3700 1498 3752 1504
rect 2504 1488 2556 1494
rect 2504 1430 2556 1436
rect 1768 1216 1820 1222
rect 1768 1158 1820 1164
rect 2228 1216 2280 1222
rect 2228 1158 2280 1164
rect 1216 1012 1268 1018
rect 1216 954 1268 960
rect 1780 950 1808 1158
rect 1847 1116 2155 1125
rect 1847 1114 1853 1116
rect 1909 1114 1933 1116
rect 1989 1114 2013 1116
rect 2069 1114 2093 1116
rect 2149 1114 2155 1116
rect 1909 1062 1911 1114
rect 2091 1062 2093 1114
rect 1847 1060 1853 1062
rect 1909 1060 1933 1062
rect 1989 1060 2013 1062
rect 2069 1060 2093 1062
rect 2149 1060 2155 1062
rect 1847 1051 2155 1060
rect 1768 944 1820 950
rect 1768 886 1820 892
rect 2240 814 2268 1158
rect 2516 1018 2544 1430
rect 2596 1420 2648 1426
rect 2596 1362 2648 1368
rect 2504 1012 2556 1018
rect 2504 954 2556 960
rect 2608 950 2636 1362
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 2813 1116 3121 1125
rect 2813 1114 2819 1116
rect 2875 1114 2899 1116
rect 2955 1114 2979 1116
rect 3035 1114 3059 1116
rect 3115 1114 3121 1116
rect 2875 1062 2877 1114
rect 3057 1062 3059 1114
rect 2813 1060 2819 1062
rect 2875 1060 2899 1062
rect 2955 1060 2979 1062
rect 3035 1060 3059 1062
rect 3115 1060 3121 1062
rect 2813 1051 3121 1060
rect 3252 1018 3280 1294
rect 3779 1116 4087 1125
rect 3779 1114 3785 1116
rect 3841 1114 3865 1116
rect 3921 1114 3945 1116
rect 4001 1114 4025 1116
rect 4081 1114 4087 1116
rect 3841 1062 3843 1114
rect 4023 1062 4025 1114
rect 3779 1060 3785 1062
rect 3841 1060 3865 1062
rect 3921 1060 3945 1062
rect 4001 1060 4025 1062
rect 4081 1060 4087 1062
rect 3779 1051 4087 1060
rect 3240 1012 3292 1018
rect 3240 954 3292 960
rect 2596 944 2648 950
rect 2596 886 2648 892
rect 664 808 716 814
rect 664 750 716 756
rect 2228 808 2280 814
rect 2228 750 2280 756
rect 3056 808 3108 814
rect 3056 750 3108 756
rect 4068 808 4120 814
rect 4068 750 4120 756
rect 676 400 704 750
rect 1860 740 1912 746
rect 1860 682 1912 688
rect 1364 572 1672 581
rect 1364 570 1370 572
rect 1426 570 1450 572
rect 1506 570 1530 572
rect 1586 570 1610 572
rect 1666 570 1672 572
rect 1426 518 1428 570
rect 1608 518 1610 570
rect 1364 516 1370 518
rect 1426 516 1450 518
rect 1506 516 1530 518
rect 1586 516 1610 518
rect 1666 516 1672 518
rect 1364 507 1672 516
rect 1872 400 1900 682
rect 2330 572 2638 581
rect 2330 570 2336 572
rect 2392 570 2416 572
rect 2472 570 2496 572
rect 2552 570 2576 572
rect 2632 570 2638 572
rect 2392 518 2394 570
rect 2574 518 2576 570
rect 2330 516 2336 518
rect 2392 516 2416 518
rect 2472 516 2496 518
rect 2552 516 2576 518
rect 2632 516 2638 518
rect 2330 507 2638 516
rect 3068 400 3096 750
rect 3296 572 3604 581
rect 3296 570 3302 572
rect 3358 570 3382 572
rect 3438 570 3462 572
rect 3518 570 3542 572
rect 3598 570 3604 572
rect 3358 518 3360 570
rect 3540 518 3542 570
rect 3296 516 3302 518
rect 3358 516 3382 518
rect 3438 516 3462 518
rect 3518 516 3542 518
rect 3598 516 3604 518
rect 3296 507 3604 516
rect 4080 474 4108 750
rect 4262 572 4570 581
rect 4262 570 4268 572
rect 4324 570 4348 572
rect 4404 570 4428 572
rect 4484 570 4508 572
rect 4564 570 4570 572
rect 4324 518 4326 570
rect 4506 518 4508 570
rect 4262 516 4268 518
rect 4324 516 4348 518
rect 4404 516 4428 518
rect 4484 516 4508 518
rect 4564 516 4570 518
rect 4262 507 4570 516
rect 4068 468 4120 474
rect 4344 468 4396 474
rect 4068 410 4120 416
rect 4264 428 4344 456
rect 4264 400 4292 428
rect 4344 410 4396 416
rect 662 0 718 400
rect 1858 0 1914 400
rect 3054 0 3110 400
rect 4250 0 4306 400
<< via2 >>
rect 887 2202 943 2204
rect 967 2202 1023 2204
rect 1047 2202 1103 2204
rect 1127 2202 1183 2204
rect 887 2150 933 2202
rect 933 2150 943 2202
rect 967 2150 997 2202
rect 997 2150 1009 2202
rect 1009 2150 1023 2202
rect 1047 2150 1061 2202
rect 1061 2150 1073 2202
rect 1073 2150 1103 2202
rect 1127 2150 1137 2202
rect 1137 2150 1183 2202
rect 887 2148 943 2150
rect 967 2148 1023 2150
rect 1047 2148 1103 2150
rect 1127 2148 1183 2150
rect 887 1114 943 1116
rect 967 1114 1023 1116
rect 1047 1114 1103 1116
rect 1127 1114 1183 1116
rect 887 1062 933 1114
rect 933 1062 943 1114
rect 967 1062 997 1114
rect 997 1062 1009 1114
rect 1009 1062 1023 1114
rect 1047 1062 1061 1114
rect 1061 1062 1073 1114
rect 1073 1062 1103 1114
rect 1127 1062 1137 1114
rect 1137 1062 1183 1114
rect 887 1060 943 1062
rect 967 1060 1023 1062
rect 1047 1060 1103 1062
rect 1127 1060 1183 1062
rect 1853 2202 1909 2204
rect 1933 2202 1989 2204
rect 2013 2202 2069 2204
rect 2093 2202 2149 2204
rect 1853 2150 1899 2202
rect 1899 2150 1909 2202
rect 1933 2150 1963 2202
rect 1963 2150 1975 2202
rect 1975 2150 1989 2202
rect 2013 2150 2027 2202
rect 2027 2150 2039 2202
rect 2039 2150 2069 2202
rect 2093 2150 2103 2202
rect 2103 2150 2149 2202
rect 1853 2148 1909 2150
rect 1933 2148 1989 2150
rect 2013 2148 2069 2150
rect 2093 2148 2149 2150
rect 2819 2202 2875 2204
rect 2899 2202 2955 2204
rect 2979 2202 3035 2204
rect 3059 2202 3115 2204
rect 2819 2150 2865 2202
rect 2865 2150 2875 2202
rect 2899 2150 2929 2202
rect 2929 2150 2941 2202
rect 2941 2150 2955 2202
rect 2979 2150 2993 2202
rect 2993 2150 3005 2202
rect 3005 2150 3035 2202
rect 3059 2150 3069 2202
rect 3069 2150 3115 2202
rect 2819 2148 2875 2150
rect 2899 2148 2955 2150
rect 2979 2148 3035 2150
rect 3059 2148 3115 2150
rect 1370 1658 1426 1660
rect 1450 1658 1506 1660
rect 1530 1658 1586 1660
rect 1610 1658 1666 1660
rect 1370 1606 1416 1658
rect 1416 1606 1426 1658
rect 1450 1606 1480 1658
rect 1480 1606 1492 1658
rect 1492 1606 1506 1658
rect 1530 1606 1544 1658
rect 1544 1606 1556 1658
rect 1556 1606 1586 1658
rect 1610 1606 1620 1658
rect 1620 1606 1666 1658
rect 1370 1604 1426 1606
rect 1450 1604 1506 1606
rect 1530 1604 1586 1606
rect 1610 1604 1666 1606
rect 2336 1658 2392 1660
rect 2416 1658 2472 1660
rect 2496 1658 2552 1660
rect 2576 1658 2632 1660
rect 2336 1606 2382 1658
rect 2382 1606 2392 1658
rect 2416 1606 2446 1658
rect 2446 1606 2458 1658
rect 2458 1606 2472 1658
rect 2496 1606 2510 1658
rect 2510 1606 2522 1658
rect 2522 1606 2552 1658
rect 2576 1606 2586 1658
rect 2586 1606 2632 1658
rect 2336 1604 2392 1606
rect 2416 1604 2472 1606
rect 2496 1604 2552 1606
rect 2576 1604 2632 1606
rect 3302 1658 3358 1660
rect 3382 1658 3438 1660
rect 3462 1658 3518 1660
rect 3542 1658 3598 1660
rect 3302 1606 3348 1658
rect 3348 1606 3358 1658
rect 3382 1606 3412 1658
rect 3412 1606 3424 1658
rect 3424 1606 3438 1658
rect 3462 1606 3476 1658
rect 3476 1606 3488 1658
rect 3488 1606 3518 1658
rect 3542 1606 3552 1658
rect 3552 1606 3598 1658
rect 3302 1604 3358 1606
rect 3382 1604 3438 1606
rect 3462 1604 3518 1606
rect 3542 1604 3598 1606
rect 3785 2202 3841 2204
rect 3865 2202 3921 2204
rect 3945 2202 4001 2204
rect 4025 2202 4081 2204
rect 3785 2150 3831 2202
rect 3831 2150 3841 2202
rect 3865 2150 3895 2202
rect 3895 2150 3907 2202
rect 3907 2150 3921 2202
rect 3945 2150 3959 2202
rect 3959 2150 3971 2202
rect 3971 2150 4001 2202
rect 4025 2150 4035 2202
rect 4035 2150 4081 2202
rect 3785 2148 3841 2150
rect 3865 2148 3921 2150
rect 3945 2148 4001 2150
rect 4025 2148 4081 2150
rect 4268 1658 4324 1660
rect 4348 1658 4404 1660
rect 4428 1658 4484 1660
rect 4508 1658 4564 1660
rect 4268 1606 4314 1658
rect 4314 1606 4324 1658
rect 4348 1606 4378 1658
rect 4378 1606 4390 1658
rect 4390 1606 4404 1658
rect 4428 1606 4442 1658
rect 4442 1606 4454 1658
rect 4454 1606 4484 1658
rect 4508 1606 4518 1658
rect 4518 1606 4564 1658
rect 4268 1604 4324 1606
rect 4348 1604 4404 1606
rect 4428 1604 4484 1606
rect 4508 1604 4564 1606
rect 1853 1114 1909 1116
rect 1933 1114 1989 1116
rect 2013 1114 2069 1116
rect 2093 1114 2149 1116
rect 1853 1062 1899 1114
rect 1899 1062 1909 1114
rect 1933 1062 1963 1114
rect 1963 1062 1975 1114
rect 1975 1062 1989 1114
rect 2013 1062 2027 1114
rect 2027 1062 2039 1114
rect 2039 1062 2069 1114
rect 2093 1062 2103 1114
rect 2103 1062 2149 1114
rect 1853 1060 1909 1062
rect 1933 1060 1989 1062
rect 2013 1060 2069 1062
rect 2093 1060 2149 1062
rect 2819 1114 2875 1116
rect 2899 1114 2955 1116
rect 2979 1114 3035 1116
rect 3059 1114 3115 1116
rect 2819 1062 2865 1114
rect 2865 1062 2875 1114
rect 2899 1062 2929 1114
rect 2929 1062 2941 1114
rect 2941 1062 2955 1114
rect 2979 1062 2993 1114
rect 2993 1062 3005 1114
rect 3005 1062 3035 1114
rect 3059 1062 3069 1114
rect 3069 1062 3115 1114
rect 2819 1060 2875 1062
rect 2899 1060 2955 1062
rect 2979 1060 3035 1062
rect 3059 1060 3115 1062
rect 3785 1114 3841 1116
rect 3865 1114 3921 1116
rect 3945 1114 4001 1116
rect 4025 1114 4081 1116
rect 3785 1062 3831 1114
rect 3831 1062 3841 1114
rect 3865 1062 3895 1114
rect 3895 1062 3907 1114
rect 3907 1062 3921 1114
rect 3945 1062 3959 1114
rect 3959 1062 3971 1114
rect 3971 1062 4001 1114
rect 4025 1062 4035 1114
rect 4035 1062 4081 1114
rect 3785 1060 3841 1062
rect 3865 1060 3921 1062
rect 3945 1060 4001 1062
rect 4025 1060 4081 1062
rect 1370 570 1426 572
rect 1450 570 1506 572
rect 1530 570 1586 572
rect 1610 570 1666 572
rect 1370 518 1416 570
rect 1416 518 1426 570
rect 1450 518 1480 570
rect 1480 518 1492 570
rect 1492 518 1506 570
rect 1530 518 1544 570
rect 1544 518 1556 570
rect 1556 518 1586 570
rect 1610 518 1620 570
rect 1620 518 1666 570
rect 1370 516 1426 518
rect 1450 516 1506 518
rect 1530 516 1586 518
rect 1610 516 1666 518
rect 2336 570 2392 572
rect 2416 570 2472 572
rect 2496 570 2552 572
rect 2576 570 2632 572
rect 2336 518 2382 570
rect 2382 518 2392 570
rect 2416 518 2446 570
rect 2446 518 2458 570
rect 2458 518 2472 570
rect 2496 518 2510 570
rect 2510 518 2522 570
rect 2522 518 2552 570
rect 2576 518 2586 570
rect 2586 518 2632 570
rect 2336 516 2392 518
rect 2416 516 2472 518
rect 2496 516 2552 518
rect 2576 516 2632 518
rect 3302 570 3358 572
rect 3382 570 3438 572
rect 3462 570 3518 572
rect 3542 570 3598 572
rect 3302 518 3348 570
rect 3348 518 3358 570
rect 3382 518 3412 570
rect 3412 518 3424 570
rect 3424 518 3438 570
rect 3462 518 3476 570
rect 3476 518 3488 570
rect 3488 518 3518 570
rect 3542 518 3552 570
rect 3552 518 3598 570
rect 3302 516 3358 518
rect 3382 516 3438 518
rect 3462 516 3518 518
rect 3542 516 3598 518
rect 4268 570 4324 572
rect 4348 570 4404 572
rect 4428 570 4484 572
rect 4508 570 4564 572
rect 4268 518 4314 570
rect 4314 518 4324 570
rect 4348 518 4378 570
rect 4378 518 4390 570
rect 4390 518 4404 570
rect 4428 518 4442 570
rect 4442 518 4454 570
rect 4454 518 4484 570
rect 4508 518 4518 570
rect 4518 518 4564 570
rect 4268 516 4324 518
rect 4348 516 4404 518
rect 4428 516 4484 518
rect 4508 516 4564 518
<< metal3 >>
rect 877 2208 1193 2209
rect 877 2144 883 2208
rect 947 2144 963 2208
rect 1027 2144 1043 2208
rect 1107 2144 1123 2208
rect 1187 2144 1193 2208
rect 877 2143 1193 2144
rect 1843 2208 2159 2209
rect 1843 2144 1849 2208
rect 1913 2144 1929 2208
rect 1993 2144 2009 2208
rect 2073 2144 2089 2208
rect 2153 2144 2159 2208
rect 1843 2143 2159 2144
rect 2809 2208 3125 2209
rect 2809 2144 2815 2208
rect 2879 2144 2895 2208
rect 2959 2144 2975 2208
rect 3039 2144 3055 2208
rect 3119 2144 3125 2208
rect 2809 2143 3125 2144
rect 3775 2208 4091 2209
rect 3775 2144 3781 2208
rect 3845 2144 3861 2208
rect 3925 2144 3941 2208
rect 4005 2144 4021 2208
rect 4085 2144 4091 2208
rect 3775 2143 4091 2144
rect 1360 1664 1676 1665
rect 1360 1600 1366 1664
rect 1430 1600 1446 1664
rect 1510 1600 1526 1664
rect 1590 1600 1606 1664
rect 1670 1600 1676 1664
rect 1360 1599 1676 1600
rect 2326 1664 2642 1665
rect 2326 1600 2332 1664
rect 2396 1600 2412 1664
rect 2476 1600 2492 1664
rect 2556 1600 2572 1664
rect 2636 1600 2642 1664
rect 2326 1599 2642 1600
rect 3292 1664 3608 1665
rect 3292 1600 3298 1664
rect 3362 1600 3378 1664
rect 3442 1600 3458 1664
rect 3522 1600 3538 1664
rect 3602 1600 3608 1664
rect 3292 1599 3608 1600
rect 4258 1664 4574 1665
rect 4258 1600 4264 1664
rect 4328 1600 4344 1664
rect 4408 1600 4424 1664
rect 4488 1600 4504 1664
rect 4568 1600 4574 1664
rect 4258 1599 4574 1600
rect 877 1120 1193 1121
rect 877 1056 883 1120
rect 947 1056 963 1120
rect 1027 1056 1043 1120
rect 1107 1056 1123 1120
rect 1187 1056 1193 1120
rect 877 1055 1193 1056
rect 1843 1120 2159 1121
rect 1843 1056 1849 1120
rect 1913 1056 1929 1120
rect 1993 1056 2009 1120
rect 2073 1056 2089 1120
rect 2153 1056 2159 1120
rect 1843 1055 2159 1056
rect 2809 1120 3125 1121
rect 2809 1056 2815 1120
rect 2879 1056 2895 1120
rect 2959 1056 2975 1120
rect 3039 1056 3055 1120
rect 3119 1056 3125 1120
rect 2809 1055 3125 1056
rect 3775 1120 4091 1121
rect 3775 1056 3781 1120
rect 3845 1056 3861 1120
rect 3925 1056 3941 1120
rect 4005 1056 4021 1120
rect 4085 1056 4091 1120
rect 3775 1055 4091 1056
rect 1360 576 1676 577
rect 1360 512 1366 576
rect 1430 512 1446 576
rect 1510 512 1526 576
rect 1590 512 1606 576
rect 1670 512 1676 576
rect 1360 511 1676 512
rect 2326 576 2642 577
rect 2326 512 2332 576
rect 2396 512 2412 576
rect 2476 512 2492 576
rect 2556 512 2572 576
rect 2636 512 2642 576
rect 2326 511 2642 512
rect 3292 576 3608 577
rect 3292 512 3298 576
rect 3362 512 3378 576
rect 3442 512 3458 576
rect 3522 512 3538 576
rect 3602 512 3608 576
rect 3292 511 3608 512
rect 4258 576 4574 577
rect 4258 512 4264 576
rect 4328 512 4344 576
rect 4408 512 4424 576
rect 4488 512 4504 576
rect 4568 512 4574 576
rect 4258 511 4574 512
<< via3 >>
rect 883 2204 947 2208
rect 883 2148 887 2204
rect 887 2148 943 2204
rect 943 2148 947 2204
rect 883 2144 947 2148
rect 963 2204 1027 2208
rect 963 2148 967 2204
rect 967 2148 1023 2204
rect 1023 2148 1027 2204
rect 963 2144 1027 2148
rect 1043 2204 1107 2208
rect 1043 2148 1047 2204
rect 1047 2148 1103 2204
rect 1103 2148 1107 2204
rect 1043 2144 1107 2148
rect 1123 2204 1187 2208
rect 1123 2148 1127 2204
rect 1127 2148 1183 2204
rect 1183 2148 1187 2204
rect 1123 2144 1187 2148
rect 1849 2204 1913 2208
rect 1849 2148 1853 2204
rect 1853 2148 1909 2204
rect 1909 2148 1913 2204
rect 1849 2144 1913 2148
rect 1929 2204 1993 2208
rect 1929 2148 1933 2204
rect 1933 2148 1989 2204
rect 1989 2148 1993 2204
rect 1929 2144 1993 2148
rect 2009 2204 2073 2208
rect 2009 2148 2013 2204
rect 2013 2148 2069 2204
rect 2069 2148 2073 2204
rect 2009 2144 2073 2148
rect 2089 2204 2153 2208
rect 2089 2148 2093 2204
rect 2093 2148 2149 2204
rect 2149 2148 2153 2204
rect 2089 2144 2153 2148
rect 2815 2204 2879 2208
rect 2815 2148 2819 2204
rect 2819 2148 2875 2204
rect 2875 2148 2879 2204
rect 2815 2144 2879 2148
rect 2895 2204 2959 2208
rect 2895 2148 2899 2204
rect 2899 2148 2955 2204
rect 2955 2148 2959 2204
rect 2895 2144 2959 2148
rect 2975 2204 3039 2208
rect 2975 2148 2979 2204
rect 2979 2148 3035 2204
rect 3035 2148 3039 2204
rect 2975 2144 3039 2148
rect 3055 2204 3119 2208
rect 3055 2148 3059 2204
rect 3059 2148 3115 2204
rect 3115 2148 3119 2204
rect 3055 2144 3119 2148
rect 3781 2204 3845 2208
rect 3781 2148 3785 2204
rect 3785 2148 3841 2204
rect 3841 2148 3845 2204
rect 3781 2144 3845 2148
rect 3861 2204 3925 2208
rect 3861 2148 3865 2204
rect 3865 2148 3921 2204
rect 3921 2148 3925 2204
rect 3861 2144 3925 2148
rect 3941 2204 4005 2208
rect 3941 2148 3945 2204
rect 3945 2148 4001 2204
rect 4001 2148 4005 2204
rect 3941 2144 4005 2148
rect 4021 2204 4085 2208
rect 4021 2148 4025 2204
rect 4025 2148 4081 2204
rect 4081 2148 4085 2204
rect 4021 2144 4085 2148
rect 1366 1660 1430 1664
rect 1366 1604 1370 1660
rect 1370 1604 1426 1660
rect 1426 1604 1430 1660
rect 1366 1600 1430 1604
rect 1446 1660 1510 1664
rect 1446 1604 1450 1660
rect 1450 1604 1506 1660
rect 1506 1604 1510 1660
rect 1446 1600 1510 1604
rect 1526 1660 1590 1664
rect 1526 1604 1530 1660
rect 1530 1604 1586 1660
rect 1586 1604 1590 1660
rect 1526 1600 1590 1604
rect 1606 1660 1670 1664
rect 1606 1604 1610 1660
rect 1610 1604 1666 1660
rect 1666 1604 1670 1660
rect 1606 1600 1670 1604
rect 2332 1660 2396 1664
rect 2332 1604 2336 1660
rect 2336 1604 2392 1660
rect 2392 1604 2396 1660
rect 2332 1600 2396 1604
rect 2412 1660 2476 1664
rect 2412 1604 2416 1660
rect 2416 1604 2472 1660
rect 2472 1604 2476 1660
rect 2412 1600 2476 1604
rect 2492 1660 2556 1664
rect 2492 1604 2496 1660
rect 2496 1604 2552 1660
rect 2552 1604 2556 1660
rect 2492 1600 2556 1604
rect 2572 1660 2636 1664
rect 2572 1604 2576 1660
rect 2576 1604 2632 1660
rect 2632 1604 2636 1660
rect 2572 1600 2636 1604
rect 3298 1660 3362 1664
rect 3298 1604 3302 1660
rect 3302 1604 3358 1660
rect 3358 1604 3362 1660
rect 3298 1600 3362 1604
rect 3378 1660 3442 1664
rect 3378 1604 3382 1660
rect 3382 1604 3438 1660
rect 3438 1604 3442 1660
rect 3378 1600 3442 1604
rect 3458 1660 3522 1664
rect 3458 1604 3462 1660
rect 3462 1604 3518 1660
rect 3518 1604 3522 1660
rect 3458 1600 3522 1604
rect 3538 1660 3602 1664
rect 3538 1604 3542 1660
rect 3542 1604 3598 1660
rect 3598 1604 3602 1660
rect 3538 1600 3602 1604
rect 4264 1660 4328 1664
rect 4264 1604 4268 1660
rect 4268 1604 4324 1660
rect 4324 1604 4328 1660
rect 4264 1600 4328 1604
rect 4344 1660 4408 1664
rect 4344 1604 4348 1660
rect 4348 1604 4404 1660
rect 4404 1604 4408 1660
rect 4344 1600 4408 1604
rect 4424 1660 4488 1664
rect 4424 1604 4428 1660
rect 4428 1604 4484 1660
rect 4484 1604 4488 1660
rect 4424 1600 4488 1604
rect 4504 1660 4568 1664
rect 4504 1604 4508 1660
rect 4508 1604 4564 1660
rect 4564 1604 4568 1660
rect 4504 1600 4568 1604
rect 883 1116 947 1120
rect 883 1060 887 1116
rect 887 1060 943 1116
rect 943 1060 947 1116
rect 883 1056 947 1060
rect 963 1116 1027 1120
rect 963 1060 967 1116
rect 967 1060 1023 1116
rect 1023 1060 1027 1116
rect 963 1056 1027 1060
rect 1043 1116 1107 1120
rect 1043 1060 1047 1116
rect 1047 1060 1103 1116
rect 1103 1060 1107 1116
rect 1043 1056 1107 1060
rect 1123 1116 1187 1120
rect 1123 1060 1127 1116
rect 1127 1060 1183 1116
rect 1183 1060 1187 1116
rect 1123 1056 1187 1060
rect 1849 1116 1913 1120
rect 1849 1060 1853 1116
rect 1853 1060 1909 1116
rect 1909 1060 1913 1116
rect 1849 1056 1913 1060
rect 1929 1116 1993 1120
rect 1929 1060 1933 1116
rect 1933 1060 1989 1116
rect 1989 1060 1993 1116
rect 1929 1056 1993 1060
rect 2009 1116 2073 1120
rect 2009 1060 2013 1116
rect 2013 1060 2069 1116
rect 2069 1060 2073 1116
rect 2009 1056 2073 1060
rect 2089 1116 2153 1120
rect 2089 1060 2093 1116
rect 2093 1060 2149 1116
rect 2149 1060 2153 1116
rect 2089 1056 2153 1060
rect 2815 1116 2879 1120
rect 2815 1060 2819 1116
rect 2819 1060 2875 1116
rect 2875 1060 2879 1116
rect 2815 1056 2879 1060
rect 2895 1116 2959 1120
rect 2895 1060 2899 1116
rect 2899 1060 2955 1116
rect 2955 1060 2959 1116
rect 2895 1056 2959 1060
rect 2975 1116 3039 1120
rect 2975 1060 2979 1116
rect 2979 1060 3035 1116
rect 3035 1060 3039 1116
rect 2975 1056 3039 1060
rect 3055 1116 3119 1120
rect 3055 1060 3059 1116
rect 3059 1060 3115 1116
rect 3115 1060 3119 1116
rect 3055 1056 3119 1060
rect 3781 1116 3845 1120
rect 3781 1060 3785 1116
rect 3785 1060 3841 1116
rect 3841 1060 3845 1116
rect 3781 1056 3845 1060
rect 3861 1116 3925 1120
rect 3861 1060 3865 1116
rect 3865 1060 3921 1116
rect 3921 1060 3925 1116
rect 3861 1056 3925 1060
rect 3941 1116 4005 1120
rect 3941 1060 3945 1116
rect 3945 1060 4001 1116
rect 4001 1060 4005 1116
rect 3941 1056 4005 1060
rect 4021 1116 4085 1120
rect 4021 1060 4025 1116
rect 4025 1060 4081 1116
rect 4081 1060 4085 1116
rect 4021 1056 4085 1060
rect 1366 572 1430 576
rect 1366 516 1370 572
rect 1370 516 1426 572
rect 1426 516 1430 572
rect 1366 512 1430 516
rect 1446 572 1510 576
rect 1446 516 1450 572
rect 1450 516 1506 572
rect 1506 516 1510 572
rect 1446 512 1510 516
rect 1526 572 1590 576
rect 1526 516 1530 572
rect 1530 516 1586 572
rect 1586 516 1590 572
rect 1526 512 1590 516
rect 1606 572 1670 576
rect 1606 516 1610 572
rect 1610 516 1666 572
rect 1666 516 1670 572
rect 1606 512 1670 516
rect 2332 572 2396 576
rect 2332 516 2336 572
rect 2336 516 2392 572
rect 2392 516 2396 572
rect 2332 512 2396 516
rect 2412 572 2476 576
rect 2412 516 2416 572
rect 2416 516 2472 572
rect 2472 516 2476 572
rect 2412 512 2476 516
rect 2492 572 2556 576
rect 2492 516 2496 572
rect 2496 516 2552 572
rect 2552 516 2556 572
rect 2492 512 2556 516
rect 2572 572 2636 576
rect 2572 516 2576 572
rect 2576 516 2632 572
rect 2632 516 2636 572
rect 2572 512 2636 516
rect 3298 572 3362 576
rect 3298 516 3302 572
rect 3302 516 3358 572
rect 3358 516 3362 572
rect 3298 512 3362 516
rect 3378 572 3442 576
rect 3378 516 3382 572
rect 3382 516 3438 572
rect 3438 516 3442 572
rect 3378 512 3442 516
rect 3458 572 3522 576
rect 3458 516 3462 572
rect 3462 516 3518 572
rect 3518 516 3522 572
rect 3458 512 3522 516
rect 3538 572 3602 576
rect 3538 516 3542 572
rect 3542 516 3598 572
rect 3598 516 3602 572
rect 3538 512 3602 516
rect 4264 572 4328 576
rect 4264 516 4268 572
rect 4268 516 4324 572
rect 4324 516 4328 572
rect 4264 512 4328 516
rect 4344 572 4408 576
rect 4344 516 4348 572
rect 4348 516 4404 572
rect 4404 516 4408 572
rect 4344 512 4408 516
rect 4424 572 4488 576
rect 4424 516 4428 572
rect 4428 516 4484 572
rect 4484 516 4488 572
rect 4424 512 4488 516
rect 4504 572 4568 576
rect 4504 516 4508 572
rect 4508 516 4564 572
rect 4564 516 4568 572
rect 4504 512 4568 516
<< metal4 >>
rect 875 2208 1195 2224
rect 875 2144 883 2208
rect 947 2144 963 2208
rect 1027 2144 1043 2208
rect 1107 2144 1123 2208
rect 1187 2144 1195 2208
rect 875 1120 1195 2144
rect 875 1056 883 1120
rect 947 1056 963 1120
rect 1027 1056 1043 1120
rect 1107 1056 1123 1120
rect 1187 1056 1195 1120
rect 875 496 1195 1056
rect 1358 1664 1678 2224
rect 1358 1600 1366 1664
rect 1430 1600 1446 1664
rect 1510 1600 1526 1664
rect 1590 1600 1606 1664
rect 1670 1600 1678 1664
rect 1358 576 1678 1600
rect 1358 512 1366 576
rect 1430 512 1446 576
rect 1510 512 1526 576
rect 1590 512 1606 576
rect 1670 512 1678 576
rect 1358 496 1678 512
rect 1841 2208 2161 2224
rect 1841 2144 1849 2208
rect 1913 2144 1929 2208
rect 1993 2144 2009 2208
rect 2073 2144 2089 2208
rect 2153 2144 2161 2208
rect 1841 1120 2161 2144
rect 1841 1056 1849 1120
rect 1913 1056 1929 1120
rect 1993 1056 2009 1120
rect 2073 1056 2089 1120
rect 2153 1056 2161 1120
rect 1841 496 2161 1056
rect 2324 1664 2644 2224
rect 2324 1600 2332 1664
rect 2396 1600 2412 1664
rect 2476 1600 2492 1664
rect 2556 1600 2572 1664
rect 2636 1600 2644 1664
rect 2324 576 2644 1600
rect 2324 512 2332 576
rect 2396 512 2412 576
rect 2476 512 2492 576
rect 2556 512 2572 576
rect 2636 512 2644 576
rect 2324 496 2644 512
rect 2807 2208 3127 2224
rect 2807 2144 2815 2208
rect 2879 2144 2895 2208
rect 2959 2144 2975 2208
rect 3039 2144 3055 2208
rect 3119 2144 3127 2208
rect 2807 1120 3127 2144
rect 2807 1056 2815 1120
rect 2879 1056 2895 1120
rect 2959 1056 2975 1120
rect 3039 1056 3055 1120
rect 3119 1056 3127 1120
rect 2807 496 3127 1056
rect 3290 1664 3610 2224
rect 3290 1600 3298 1664
rect 3362 1600 3378 1664
rect 3442 1600 3458 1664
rect 3522 1600 3538 1664
rect 3602 1600 3610 1664
rect 3290 576 3610 1600
rect 3290 512 3298 576
rect 3362 512 3378 576
rect 3442 512 3458 576
rect 3522 512 3538 576
rect 3602 512 3610 576
rect 3290 496 3610 512
rect 3773 2208 4093 2224
rect 3773 2144 3781 2208
rect 3845 2144 3861 2208
rect 3925 2144 3941 2208
rect 4005 2144 4021 2208
rect 4085 2144 4093 2208
rect 3773 1120 4093 2144
rect 3773 1056 3781 1120
rect 3845 1056 3861 1120
rect 3925 1056 3941 1120
rect 4005 1056 4021 1120
rect 4085 1056 4093 1120
rect 3773 496 4093 1056
rect 4256 1664 4576 2224
rect 4256 1600 4264 1664
rect 4328 1600 4344 1664
rect 4408 1600 4424 1664
rect 4488 1600 4504 1664
rect 4568 1600 4576 1664
rect 4256 576 4576 1600
rect 4256 512 4264 576
rect 4328 512 4344 576
rect 4408 512 4424 576
rect 4488 512 4504 576
rect 4568 512 4576 576
rect 4256 496 4576 512
use sky130_fd_sc_hd__xnor2_1  _3_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2852 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _4_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1748 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _5_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2300 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _6_
timestamp 1704896540
transform 1 0 2852 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _7_
timestamp 1704896540
transform 1 0 3312 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1104 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1840 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2576 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3496 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1564 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_34
timestamp 1704896540
transform 1 0 3680 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_38
timestamp 1704896540
transform 1 0 4048 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3220 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_37
timestamp 1704896540
transform 1 0 3956 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 1104 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1704896540
transform -1 0 2576 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform 1 0 3864 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 4416 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_4
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 4416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_5
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 4416 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_7
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
<< labels >>
rlabel metal2 s 2564 1632 2564 1632 4 VGND
rlabel metal1 s 2484 2176 2484 2176 4 VPWR
rlabel metal1 s 3312 1394 3312 1394 4 _0_
rlabel metal1 s 2129 1530 2129 1530 4 _1_
rlabel metal2 s 2254 986 2254 986 4 _2_
rlabel metal2 s 690 568 690 568 4 analog_to_digital_in[0]
rlabel metal2 s 1886 534 1886 534 4 analog_to_digital_in[1]
rlabel metal2 s 3082 568 3082 568 4 analog_to_digital_in[2]
rlabel metal2 s 4250 0 4306 400 4 analog_to_digital_in[3]
port 6 nsew
rlabel metal1 s 1656 986 1656 986 4 encoded_out[0]
rlabel metal1 s 3634 1530 3634 1530 4 encoded_out[1]
rlabel metal1 s 1886 1190 1886 1190 4 net1
rlabel metal1 s 2346 1462 2346 1462 4 net2
rlabel metal1 s 2990 1326 2990 1326 4 net3
rlabel metal1 s 3266 918 3266 918 4 net4
flabel metal4 s 4256 496 4576 2224 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3290 496 3610 2224 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2324 496 2644 2224 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 1358 496 1678 2224 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 3773 496 4093 2224 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2807 496 3127 2224 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1841 496 2161 2224 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 875 496 1195 2224 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 662 0 718 400 0 FreeSans 280 90 0 0 analog_to_digital_in[0]
port 3 nsew
flabel metal2 s 1858 0 1914 400 0 FreeSans 280 90 0 0 analog_to_digital_in[1]
port 4 nsew
flabel metal2 s 3054 0 3110 400 0 FreeSans 280 90 0 0 analog_to_digital_in[2]
port 5 nsew
flabel metal2 s 4278 200 4278 200 0 FreeSans 280 90 0 0 analog_to_digital_in[3]
flabel metal2 s 1214 2600 1270 3000 0 FreeSans 280 90 0 0 encoded_out[0]
port 7 nsew
flabel metal2 s 3698 2600 3754 3000 0 FreeSans 280 90 0 0 encoded_out[1]
port 8 nsew
<< properties >>
string FIXED_BBOX 0 0 5000 3000
string GDS_END 74508
string GDS_FILE ../gds/adc_digital_control.gds
string GDS_START 41232
<< end >>
