** sch_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp_ladder.sch
.subckt opamp_ladder VDD in VSS out3 out2 out1 out0
*.PININFO out0:O out2:O out3:O in:I VDD:B VSS:B out1:O
x1 VDD node_0 in out0 VSS opamp
x2 VDD node_1 in out1 VSS opamp
x3 VDD node_2 in out2 VSS opamp
x4 VDD node_3 in out3 VSS opamp
XR1 node_3 VDD VSS sky130_fd_pr__res_high_po_0p69 L=7.34 mult=1 m=1
XR2 node_2 node_3 VSS sky130_fd_pr__res_high_po_0p69 L=3.45 mult=1 m=1
XR3 node_1 node_2 VSS sky130_fd_pr__res_high_po_0p69 L=3.45 mult=1 m=1
XR4 node_0 node_1 VSS sky130_fd_pr__res_high_po_0p69 L=3.45 mult=1 m=1
XR5 VSS node_0 VSS sky130_fd_pr__res_high_po_0p69 L=3.45 mult=1 m=1
.ends

* expanding   symbol:  opamp.sym # of pins=5
** sym_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp.sym
** sch_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp.sch
.subckt opamp VDD vin_n vin_p Vout VGND
*.PININFO vin_n:I vin_p:I Vout:O VDD:B VGND:B
XM1 net1 vin_n net3 VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 m=1
XM2 net2 vin_p net3 VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 m=1
XM3 net1 net1 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 m=1
XM4 net2 net1 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 m=1
XM5 net3 net4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 m=1
XM7 Vout net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 m=1
XM8 net4 net4 VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 m=1
XM6 Vout net2 VGND VGND sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 m=1
XR VGND net8 VGND sky130_fd_pr__res_high_po_0p35 L=4 mult=1 m=1
XR1 net8 net7 VGND sky130_fd_pr__res_high_po_0p35 L=4 mult=1 m=1
XR2 net7 net6 VGND sky130_fd_pr__res_high_po_0p35 L=4 mult=1 m=1
XR3 net6 net5 VGND sky130_fd_pr__res_high_po_0p35 L=4 mult=1 m=1
XR4 net5 net4 VGND sky130_fd_pr__res_high_po_0p35 L=4 mult=1 m=1
.ends

.end
