** sch_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp_ladder_tb.sch
**.subckt opamp_ladder_tb out0 out1 out2 out3 in
*.opin out0
*.opin out1
*.opin out2
*.opin out3
*.ipin in
x1 VDD in VSS out3 out2 out1 out0 opamp_ladder
V1 VSS GND 0
V2 VDD GND 1.8
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ttuser/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt





v_in in 0 1.8
.control
dc v_in 0 1.8 0.01
save all
write opamp_ladder_tb.raw
.endc



**** end user architecture code
**.ends

* expanding   symbol:  opamp_ladder.sym # of pins=7
** sym_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp_ladder.sym
** sch_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp_ladder.sch
.subckt opamp_ladder VDD in VSS out3 out2 out1 out0
*.opin out0
*.opin out2
*.opin out3
*.ipin in
*.iopin VDD
*.iopin VSS
*.opin out1
x1 VDD VSS net4 in out0 VSS opamp
XR2 VSS net4 VSS sky130_fd_pr__res_generic_nd W=1 L=8.4 mult=1 m=1
XR3 net4 net3 VSS sky130_fd_pr__res_generic_nd W=1 L=8.4 mult=1 m=1
XR4 net3 net2 VSS sky130_fd_pr__res_generic_nd W=1 L=8.4 mult=1 m=1
XR5 net2 net1 VSS sky130_fd_pr__res_generic_nd W=1 L=8.4 mult=1 m=1
x2 VDD VSS net3 in out1 VSS opamp
x3 VDD VSS net2 in out2 VSS opamp
x4 VDD VSS net1 in out3 VSS opamp
XR1 net1 VDD VSS sky130_fd_pr__res_generic_nd W=1 L=8.4 mult=1 m=1
.ends


* expanding   symbol:  opamp.sym # of pins=6
** sym_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp.sym
** sch_path: /home/ttuser/Documents/tt08-analog-adc/xschem/opamp.sch
.subckt opamp VDD ZREF vin_n vin_p Vout VGND
*.ipin vin_n
*.ipin vin_p
*.opin Vout
*.iopin VDD
*.iopin ZREF
*.iopin VGND
XM1 net1 vin_n net3 net3 sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 vin_p net3 net3 sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 net1 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 net1 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net3 VGND VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vout VGND VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 ZREF VGND VDD VDD sky130_fd_pr__pfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net4 VDD net2 VGND sky130_fd_pr__nfet_01v8 L=0.6 W=1 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)' nrd='0.29 / W'
+ nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XC1 net4 Vout sky130_fd_pr__cap_mim_m3_1 W=17.55 L=15 MF=1 m=1
XM6 Vout net2 VGND VGND sky130_fd_pr__nfet_01v8 L=0.6 W=6 nf=1 ad='W * 0.29' as='W * 0.29' pd='2 * (W + 0.29)' ps='2 * (W + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XR1 ZREF VDD VGND sky130_fd_pr__res_generic_nd W=1 L=5 mult=1 m=1
XR2 VGND ZREF VGND sky130_fd_pr__res_generic_nd W=1 L=5 mult=1 m=1
.ends

.GLOBAL GND
.end
