magic
tech sky130A
timestamp 1728463006
<< error_p >>
rect 17636 7850 17664 7864
rect 17636 7836 17650 7850
rect 17636 7775 17664 7789
rect 17711 7775 17764 7789
rect 17650 7764 17675 7775
rect 17725 7764 17750 7775
rect 17650 7750 17689 7764
rect 17675 7736 17689 7750
rect 17711 7750 17750 7764
rect 17711 7736 17725 7750
rect 9422 7497 9475 7500
rect 5350 7100 5375 7103
rect 5350 7072 5375 7075
rect 5350 7025 5375 7028
rect 5350 6997 5375 7000
rect 5350 6950 5375 6953
rect 5350 6922 5375 6925
rect 5350 6900 5375 6903
rect 5350 6872 5375 6875
rect 5350 6822 5375 6825
rect 5350 6772 5375 6775
<< metal2 >>
rect 15150 8425 16000 8450
rect 14975 8400 16175 8425
rect 14875 8375 16325 8400
rect 14800 8350 16425 8375
rect 14750 8325 16525 8350
rect 14725 8300 16625 8325
rect 4675 7600 5175 8300
rect 9250 8275 9400 8300
rect 11450 8275 11700 8300
rect 14700 8275 16700 8300
rect 9225 8250 9425 8275
rect 11450 8250 11725 8275
rect 14650 8250 16750 8275
rect 9225 8225 9450 8250
rect 11450 8225 11750 8250
rect 14550 8225 16825 8250
rect 9200 8200 9475 8225
rect 11450 8200 11775 8225
rect 14500 8200 16875 8225
rect 9175 8175 9500 8200
rect 9150 8150 9525 8175
rect 9125 8125 9525 8150
rect 11450 8150 11800 8200
rect 14425 8175 15325 8200
rect 15625 8175 16925 8200
rect 14375 8150 15050 8175
rect 15875 8150 16975 8175
rect 11450 8125 11825 8150
rect 14300 8125 14900 8150
rect 16025 8125 17025 8150
rect 9100 8100 9550 8125
rect 11450 8100 11850 8125
rect 14250 8100 14800 8125
rect 16125 8100 17050 8125
rect 9075 8075 9575 8100
rect 11450 8075 11875 8100
rect 14200 8075 14700 8100
rect 16225 8075 17100 8100
rect 9050 8050 9600 8075
rect 11450 8050 11900 8075
rect 14175 8050 14600 8075
rect 16300 8050 17125 8075
rect 6625 8025 6650 8050
rect 9025 8025 9625 8050
rect 11450 8025 11925 8050
rect 14125 8025 14550 8050
rect 16375 8025 17150 8050
rect 6625 8000 6875 8025
rect 9000 8000 9650 8025
rect 11450 8000 11950 8025
rect 14100 8000 14475 8025
rect 16425 8000 17200 8025
rect 6625 7975 6950 8000
rect 8975 7975 9675 8000
rect 11450 7975 11975 8000
rect 14050 7975 14425 8000
rect 16500 7975 17225 8000
rect 6625 7950 7000 7975
rect 8975 7950 9700 7975
rect 6625 7925 7025 7950
rect 8950 7925 9725 7950
rect 11450 7925 12000 7975
rect 14025 7950 14375 7975
rect 16550 7950 17250 7975
rect 14000 7925 14325 7950
rect 16600 7925 17275 7950
rect 6625 7900 7075 7925
rect 8925 7900 9750 7925
rect 6625 7850 7100 7900
rect 8900 7875 9750 7900
rect 11450 7900 12025 7925
rect 13975 7900 14275 7925
rect 16625 7900 17300 7925
rect 8875 7850 9100 7875
rect 9150 7850 9775 7875
rect 6625 7825 7125 7850
rect 8850 7825 9075 7850
rect 9175 7825 9800 7850
rect 6625 7775 7150 7825
rect 8825 7800 9050 7825
rect 9200 7800 9825 7825
rect 8800 7775 9025 7800
rect 9225 7775 9850 7800
rect 4675 7575 5200 7600
rect 4675 7550 5225 7575
rect 4675 7525 5250 7550
rect 6625 7525 7175 7775
rect 9250 7750 9875 7775
rect 9275 7725 9900 7750
rect 9275 7700 9925 7725
rect 9300 7675 9950 7700
rect 9325 7650 9975 7675
rect 9350 7625 10000 7650
rect 9375 7600 10000 7625
rect 9400 7575 10025 7600
rect 9425 7550 10050 7575
rect 9450 7525 10075 7550
rect 4675 7325 7175 7525
rect 9475 7500 10100 7525
rect 8550 7475 10125 7500
rect 8525 7450 10150 7475
rect 8500 7425 10175 7450
rect 8475 7400 10200 7425
rect 8450 7375 10225 7400
rect 8425 7350 10225 7375
rect 8400 7325 10250 7350
rect 4675 7125 5350 7325
rect 4675 7100 5375 7125
rect 4675 7075 5350 7100
rect 4675 7025 5375 7075
rect 4675 7000 5350 7025
rect 4675 6950 5375 7000
rect 4675 6925 5350 6950
rect 4675 6900 5375 6925
rect 4675 6875 5350 6900
rect 4675 6850 5375 6875
rect 4675 6825 5350 6850
rect 4675 6800 5375 6825
rect 4675 6775 5350 6800
rect 4675 6750 5375 6775
rect 4675 6575 5350 6750
rect 6625 6625 7175 7325
rect 8375 7300 10275 7325
rect 8350 7275 8975 7300
rect 9650 7275 10300 7300
rect 8325 7250 8925 7275
rect 9675 7250 10325 7275
rect 8325 7225 8900 7250
rect 9700 7225 10350 7250
rect 8300 7200 8875 7225
rect 9725 7200 10375 7225
rect 8275 7175 8850 7200
rect 9725 7175 10400 7200
rect 8250 7150 8825 7175
rect 9750 7150 10425 7175
rect 8225 7125 8800 7150
rect 9775 7125 10450 7150
rect 8200 7100 8800 7125
rect 9800 7100 10450 7125
rect 8175 7075 8775 7100
rect 9825 7075 10475 7100
rect 8150 7050 8750 7075
rect 9850 7050 10500 7075
rect 8125 7025 8725 7050
rect 9875 7025 10525 7050
rect 8100 7000 8700 7025
rect 9900 7000 10550 7025
rect 11450 7000 12050 7900
rect 13950 7875 14250 7900
rect 16675 7875 17325 7900
rect 13925 7850 14200 7875
rect 16700 7850 17350 7875
rect 17650 7850 17750 7875
rect 13900 7825 14175 7850
rect 16750 7825 17350 7850
rect 13900 7800 14150 7825
rect 16775 7800 17375 7825
rect 13875 7775 14125 7800
rect 16800 7775 17400 7800
rect 17625 7775 17650 7850
rect 17675 7800 17725 7850
rect 17700 7775 17725 7800
rect 17750 7775 17775 7825
rect 13850 7750 14100 7775
rect 16825 7750 17400 7775
rect 17650 7750 17675 7775
rect 17725 7750 17750 7775
rect 13875 7725 14075 7750
rect 16850 7725 17425 7750
rect 17675 7725 17725 7750
rect 13950 7700 14050 7725
rect 14025 7675 14050 7700
rect 16875 7700 17425 7725
rect 16875 7675 17450 7700
rect 15400 7650 15600 7675
rect 16900 7650 17450 7675
rect 15300 7625 15700 7650
rect 16900 7625 17475 7650
rect 15250 7600 15750 7625
rect 16900 7600 17550 7625
rect 17575 7600 17625 7625
rect 17775 7600 17800 7625
rect 15225 7575 15775 7600
rect 15200 7550 15800 7575
rect 15200 7525 15825 7550
rect 15175 7475 15825 7525
rect 16925 7475 17825 7600
rect 15200 7425 15800 7475
rect 16900 7450 17500 7475
rect 16900 7425 17475 7450
rect 15225 7400 15775 7425
rect 15275 7375 15725 7400
rect 16875 7375 17450 7425
rect 15325 7350 15675 7375
rect 16850 7350 17425 7375
rect 15475 7325 15525 7350
rect 16825 7325 17425 7350
rect 16825 7300 17400 7325
rect 16800 7275 17375 7300
rect 16750 7250 17375 7275
rect 16725 7225 17350 7250
rect 16700 7200 17325 7225
rect 16650 7175 17300 7200
rect 16625 7150 17275 7175
rect 16575 7125 17250 7150
rect 16525 7100 17225 7125
rect 16475 7075 17200 7100
rect 16400 7050 17175 7075
rect 16350 7025 17150 7050
rect 14625 7000 14650 7025
rect 16275 7000 17125 7025
rect 8075 6975 8675 7000
rect 9925 6975 10575 7000
rect 8075 6950 8650 6975
rect 9950 6950 10600 6975
rect 11450 6950 12075 7000
rect 14625 6975 14725 7000
rect 16175 6975 17075 7000
rect 14600 6950 14850 6975
rect 16075 6950 17050 6975
rect 8050 6925 8625 6950
rect 9975 6925 10625 6950
rect 11450 6925 12100 6950
rect 14575 6925 14975 6950
rect 15950 6925 17000 6950
rect 8025 6900 8600 6925
rect 10000 6900 10650 6925
rect 11450 6900 12125 6925
rect 14575 6900 15150 6925
rect 15775 6900 16950 6925
rect 8000 6875 8575 6900
rect 7975 6850 8550 6875
rect 10025 6850 10675 6900
rect 11450 6875 12225 6900
rect 14550 6875 16900 6900
rect 11450 6850 13525 6875
rect 14550 6850 16850 6875
rect 7950 6825 8550 6850
rect 10050 6825 10700 6850
rect 11475 6825 13550 6850
rect 14575 6825 16800 6850
rect 7925 6800 8525 6825
rect 10075 6800 10725 6825
rect 11500 6800 13575 6825
rect 14650 6800 16750 6825
rect 7900 6775 8500 6800
rect 10100 6775 10750 6800
rect 11525 6775 13600 6800
rect 14750 6775 16675 6800
rect 7875 6750 8475 6775
rect 10125 6750 10775 6775
rect 11550 6750 13650 6775
rect 14850 6750 16600 6775
rect 7850 6725 8450 6750
rect 10150 6725 10800 6750
rect 11575 6725 13675 6750
rect 15000 6725 16500 6750
rect 7850 6700 8425 6725
rect 10175 6700 10825 6725
rect 11575 6700 13700 6725
rect 15225 6700 16400 6725
rect 7825 6675 8400 6700
rect 10200 6675 10850 6700
rect 11600 6675 13700 6700
rect 15275 6675 16275 6700
rect 7800 6650 8375 6675
rect 10225 6650 10875 6675
rect 11625 6650 13700 6675
rect 15300 6650 16100 6675
rect 7775 6625 8350 6650
rect 10250 6625 10900 6650
rect 11650 6625 13700 6650
rect 15325 6625 15875 6650
rect 10275 6600 10900 6625
rect 4675 6550 5375 6575
<< end >>
